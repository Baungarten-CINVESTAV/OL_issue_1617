magic
tech sky130A
magscale 1 2
timestamp 1674174216
<< viali >>
rect 14473 37417 14507 37451
rect 26525 37417 26559 37451
rect 32505 37417 32539 37451
rect 34253 37417 34287 37451
rect 5917 37281 5951 37315
rect 6745 37281 6779 37315
rect 7481 37281 7515 37315
rect 27169 37281 27203 37315
rect 32965 37281 32999 37315
rect 34897 37281 34931 37315
rect 2329 37213 2363 37247
rect 3065 37213 3099 37247
rect 4261 37213 4295 37247
rect 5457 37213 5491 37247
rect 7297 37213 7331 37247
rect 9413 37213 9447 37247
rect 10701 37213 10735 37247
rect 11713 37213 11747 37247
rect 13737 37213 13771 37247
rect 15117 37213 15151 37247
rect 16865 37213 16899 37247
rect 18337 37213 18371 37247
rect 18797 37213 18831 37247
rect 20085 37213 20119 37247
rect 22017 37213 22051 37247
rect 22845 37213 22879 37247
rect 23305 37213 23339 37247
rect 24593 37213 24627 37247
rect 27445 37213 27479 37247
rect 28457 37213 28491 37247
rect 29745 37213 29779 37247
rect 31033 37213 31067 37247
rect 33149 37213 33183 37247
rect 35081 37213 35115 37247
rect 36093 37213 36127 37247
rect 2145 37077 2179 37111
rect 2881 37077 2915 37111
rect 4077 37077 4111 37111
rect 5273 37077 5307 37111
rect 9229 37077 9263 37111
rect 10517 37077 10551 37111
rect 11897 37077 11931 37111
rect 13553 37077 13587 37111
rect 15025 37077 15059 37111
rect 17049 37077 17083 37111
rect 18153 37077 18187 37111
rect 20269 37077 20303 37111
rect 22201 37077 22235 37111
rect 23489 37077 23523 37111
rect 24777 37077 24811 37111
rect 28641 37077 28675 37111
rect 29929 37077 29963 37111
rect 31217 37077 31251 37111
rect 36277 37077 36311 37111
rect 11713 36873 11747 36907
rect 27353 36873 27387 36907
rect 29101 36873 29135 36907
rect 31309 36873 31343 36907
rect 35541 36873 35575 36907
rect 1685 36805 1719 36839
rect 2329 36805 2363 36839
rect 34897 36805 34931 36839
rect 36277 36805 36311 36839
rect 11897 36737 11931 36771
rect 27169 36737 27203 36771
rect 27813 36737 27847 36771
rect 28917 36737 28951 36771
rect 31125 36737 31159 36771
rect 35357 36737 35391 36771
rect 1869 36601 1903 36635
rect 3249 36533 3283 36567
rect 13921 36533 13955 36567
rect 28365 36533 28399 36567
rect 36185 36533 36219 36567
rect 35633 36329 35667 36363
rect 1777 36261 1811 36295
rect 26709 36261 26743 36295
rect 1593 36125 1627 36159
rect 2237 36125 2271 36159
rect 26525 36125 26559 36159
rect 27169 36125 27203 36159
rect 36093 36125 36127 36159
rect 36277 35989 36311 36023
rect 1593 35581 1627 35615
rect 1869 35581 1903 35615
rect 1593 35241 1627 35275
rect 36093 35037 36127 35071
rect 36369 35037 36403 35071
rect 36369 34697 36403 34731
rect 18889 33065 18923 33099
rect 18705 32861 18739 32895
rect 19441 32861 19475 32895
rect 24593 32861 24627 32895
rect 25237 32861 25271 32895
rect 24685 32793 24719 32827
rect 35633 32793 35667 32827
rect 36277 32793 36311 32827
rect 36185 32725 36219 32759
rect 1593 32317 1627 32351
rect 1869 32317 1903 32351
rect 1593 31977 1627 32011
rect 10057 31977 10091 32011
rect 36277 31909 36311 31943
rect 9965 31773 9999 31807
rect 10701 31773 10735 31807
rect 10793 31773 10827 31807
rect 36093 31773 36127 31807
rect 10333 31433 10367 31467
rect 10425 31297 10459 31331
rect 21373 30889 21407 30923
rect 1869 30685 1903 30719
rect 21281 30685 21315 30719
rect 1685 30549 1719 30583
rect 13185 30345 13219 30379
rect 4905 30277 4939 30311
rect 4813 30209 4847 30243
rect 12449 30209 12483 30243
rect 13369 30209 13403 30243
rect 22661 30209 22695 30243
rect 12265 30073 12299 30107
rect 13921 30073 13955 30107
rect 22569 30005 22603 30039
rect 22201 29597 22235 29631
rect 22753 29597 22787 29631
rect 35633 29529 35667 29563
rect 36277 29529 36311 29563
rect 12541 29461 12575 29495
rect 22109 29461 22143 29495
rect 36185 29461 36219 29495
rect 16129 29257 16163 29291
rect 1593 29121 1627 29155
rect 2237 29121 2271 29155
rect 15669 29121 15703 29155
rect 1777 28985 1811 29019
rect 15577 28985 15611 29019
rect 14657 28713 14691 28747
rect 14473 28509 14507 28543
rect 15117 28509 15151 28543
rect 35633 28033 35667 28067
rect 36277 28033 36311 28067
rect 15301 27897 15335 27931
rect 36093 27897 36127 27931
rect 1961 27829 1995 27863
rect 11989 27829 12023 27863
rect 15761 27829 15795 27863
rect 12633 27557 12667 27591
rect 1869 27421 1903 27455
rect 2513 27421 2547 27455
rect 15577 27421 15611 27455
rect 16037 27353 16071 27387
rect 1685 27285 1719 27319
rect 2329 27285 2363 27319
rect 10885 27285 10919 27319
rect 11713 27285 11747 27319
rect 14381 27285 14415 27319
rect 14841 27285 14875 27319
rect 15485 27285 15519 27319
rect 8033 27013 8067 27047
rect 11805 27013 11839 27047
rect 11897 27013 11931 27047
rect 13093 27013 13127 27047
rect 13645 27013 13679 27047
rect 14933 27013 14967 27047
rect 15025 27013 15059 27047
rect 15669 27013 15703 27047
rect 15761 27013 15795 27047
rect 2145 26945 2179 26979
rect 2789 26945 2823 26979
rect 11161 26945 11195 26979
rect 17049 26945 17083 26979
rect 17509 26945 17543 26979
rect 7941 26877 7975 26911
rect 12449 26877 12483 26911
rect 13001 26877 13035 26911
rect 14749 26877 14783 26911
rect 16313 26877 16347 26911
rect 2605 26809 2639 26843
rect 8493 26809 8527 26843
rect 2053 26741 2087 26775
rect 10517 26741 10551 26775
rect 11069 26741 11103 26775
rect 16957 26741 16991 26775
rect 11713 26537 11747 26571
rect 1685 26469 1719 26503
rect 10517 26469 10551 26503
rect 12357 26469 12391 26503
rect 36277 26469 36311 26503
rect 2421 26401 2455 26435
rect 7941 26401 7975 26435
rect 9229 26401 9263 26435
rect 9873 26401 9907 26435
rect 11069 26401 11103 26435
rect 12909 26401 12943 26435
rect 13553 26401 13587 26435
rect 16037 26401 16071 26435
rect 16681 26401 16715 26435
rect 17325 26401 17359 26435
rect 18797 26401 18831 26435
rect 1869 26333 1903 26367
rect 2513 26333 2547 26367
rect 11621 26333 11655 26367
rect 12449 26333 12483 26367
rect 14933 26333 14967 26367
rect 36093 26333 36127 26367
rect 2973 26265 3007 26299
rect 9781 26265 9815 26299
rect 10977 26265 11011 26299
rect 13461 26265 13495 26299
rect 15393 26265 15427 26299
rect 15945 26265 15979 26299
rect 16773 26265 16807 26299
rect 18153 26265 18187 26299
rect 18705 26265 18739 26299
rect 14841 26197 14875 26231
rect 8585 25993 8619 26027
rect 9321 25993 9355 26027
rect 2145 25925 2179 25959
rect 5273 25925 5307 25959
rect 13277 25925 13311 25959
rect 14381 25925 14415 25959
rect 14933 25925 14967 25959
rect 17417 25925 17451 25959
rect 2789 25857 2823 25891
rect 3433 25857 3467 25891
rect 8677 25857 8711 25891
rect 9229 25857 9263 25891
rect 9873 25857 9907 25891
rect 10977 25857 11011 25891
rect 12081 25857 12115 25891
rect 15577 25857 15611 25891
rect 16037 25857 16071 25891
rect 18245 25857 18279 25891
rect 18797 25857 18831 25891
rect 1961 25789 1995 25823
rect 2237 25789 2271 25823
rect 5181 25789 5215 25823
rect 7205 25789 7239 25823
rect 12725 25789 12759 25823
rect 13369 25789 13403 25823
rect 14289 25789 14323 25823
rect 17509 25789 17543 25823
rect 2881 25721 2915 25755
rect 5733 25721 5767 25755
rect 16957 25721 16991 25755
rect 3525 25653 3559 25687
rect 7941 25653 7975 25687
rect 9965 25653 9999 25687
rect 11069 25653 11103 25687
rect 12173 25653 12207 25687
rect 15485 25653 15519 25687
rect 16129 25653 16163 25687
rect 18153 25653 18187 25687
rect 17049 25449 17083 25483
rect 6285 25381 6319 25415
rect 18245 25381 18279 25415
rect 20361 25381 20395 25415
rect 2237 25313 2271 25347
rect 4077 25313 4111 25347
rect 10977 25313 11011 25347
rect 11345 25313 11379 25347
rect 12265 25313 12299 25347
rect 14289 25313 14323 25347
rect 17693 25313 17727 25347
rect 20913 25313 20947 25347
rect 3341 25245 3375 25279
rect 4629 25245 4663 25279
rect 9321 25245 9355 25279
rect 9965 25245 9999 25279
rect 12081 25245 12115 25279
rect 13553 25245 13587 25279
rect 13645 25245 13679 25279
rect 15209 25245 15243 25279
rect 15945 25245 15979 25279
rect 16957 25245 16991 25279
rect 2421 25177 2455 25211
rect 2513 25177 2547 25211
rect 5733 25177 5767 25211
rect 5825 25177 5859 25211
rect 6929 25177 6963 25211
rect 7021 25177 7055 25211
rect 7573 25177 7607 25211
rect 8585 25177 8619 25211
rect 11253 25177 11287 25211
rect 12725 25177 12759 25211
rect 14473 25177 14507 25211
rect 17785 25177 17819 25211
rect 20821 25177 20855 25211
rect 3157 25109 3191 25143
rect 5181 25109 5215 25143
rect 9873 25109 9907 25143
rect 15301 25109 15335 25143
rect 16037 25109 16071 25143
rect 18797 25109 18831 25143
rect 19441 25109 19475 25143
rect 2145 24837 2179 24871
rect 3893 24837 3927 24871
rect 10517 24837 10551 24871
rect 11897 24837 11931 24871
rect 13645 24837 13679 24871
rect 14841 24837 14875 24871
rect 17049 24837 17083 24871
rect 2789 24769 2823 24803
rect 5825 24769 5859 24803
rect 5917 24769 5951 24803
rect 6561 24769 6595 24803
rect 7389 24769 7423 24803
rect 8033 24769 8067 24803
rect 8677 24769 8711 24803
rect 9413 24769 9447 24803
rect 9505 24769 9539 24803
rect 14197 24769 14231 24803
rect 18521 24769 18555 24803
rect 18613 24769 18647 24803
rect 2237 24701 2271 24735
rect 3709 24701 3743 24735
rect 3985 24701 4019 24735
rect 6653 24701 6687 24735
rect 7481 24701 7515 24735
rect 10609 24701 10643 24735
rect 11805 24701 11839 24735
rect 13553 24701 13587 24735
rect 14749 24701 14783 24735
rect 15761 24701 15795 24735
rect 16957 24701 16991 24735
rect 17233 24701 17267 24735
rect 19073 24701 19107 24735
rect 36093 24701 36127 24735
rect 36369 24701 36403 24735
rect 1685 24633 1719 24667
rect 5365 24633 5399 24667
rect 8769 24633 8803 24667
rect 10057 24633 10091 24667
rect 12357 24633 12391 24667
rect 4629 24565 4663 24599
rect 8125 24565 8159 24599
rect 13001 24565 13035 24599
rect 16313 24565 16347 24599
rect 19717 24565 19751 24599
rect 2237 24361 2271 24395
rect 3985 24361 4019 24395
rect 6377 24361 6411 24395
rect 7021 24361 7055 24395
rect 20913 24361 20947 24395
rect 36369 24361 36403 24395
rect 10057 24293 10091 24327
rect 2881 24225 2915 24259
rect 8493 24225 8527 24259
rect 9505 24225 9539 24259
rect 10701 24225 10735 24259
rect 11345 24225 11379 24259
rect 12173 24225 12207 24259
rect 12449 24225 12483 24259
rect 13093 24225 13127 24259
rect 13369 24225 13403 24259
rect 14657 24225 14691 24259
rect 15577 24225 15611 24259
rect 16681 24225 16715 24259
rect 17969 24225 18003 24259
rect 18245 24225 18279 24259
rect 2329 24157 2363 24191
rect 2789 24157 2823 24191
rect 4169 24157 4203 24191
rect 5181 24157 5215 24191
rect 6469 24157 6503 24191
rect 7113 24157 7147 24191
rect 7757 24157 7791 24191
rect 7849 24157 7883 24191
rect 8401 24157 8435 24191
rect 17417 24157 17451 24191
rect 19901 24157 19935 24191
rect 21005 24157 21039 24191
rect 5273 24089 5307 24123
rect 9597 24089 9631 24123
rect 10793 24089 10827 24123
rect 12357 24089 12391 24123
rect 13185 24089 13219 24123
rect 14381 24089 14415 24123
rect 14473 24089 14507 24123
rect 16037 24089 16071 24123
rect 16589 24089 16623 24123
rect 18061 24089 18095 24123
rect 1593 24021 1627 24055
rect 4629 24021 4663 24055
rect 17325 24021 17359 24055
rect 19993 24021 20027 24055
rect 21465 24021 21499 24055
rect 14013 23817 14047 23851
rect 27813 23817 27847 23851
rect 5457 23749 5491 23783
rect 8125 23749 8159 23783
rect 8217 23749 8251 23783
rect 8953 23749 8987 23783
rect 9505 23749 9539 23783
rect 10977 23749 11011 23783
rect 11069 23749 11103 23783
rect 12725 23749 12759 23783
rect 12817 23749 12851 23783
rect 16129 23749 16163 23783
rect 17049 23749 17083 23783
rect 17601 23749 17635 23783
rect 19717 23749 19751 23783
rect 20269 23749 20303 23783
rect 2237 23681 2271 23715
rect 2697 23681 2731 23715
rect 2789 23681 2823 23715
rect 3525 23681 3559 23715
rect 3985 23681 4019 23715
rect 6929 23681 6963 23715
rect 12173 23681 12207 23715
rect 13369 23681 13403 23715
rect 19073 23681 19107 23715
rect 22201 23681 22235 23715
rect 27629 23681 27663 23715
rect 28273 23681 28307 23715
rect 5365 23613 5399 23647
rect 5733 23613 5767 23647
rect 7573 23613 7607 23647
rect 8861 23613 8895 23647
rect 10793 23613 10827 23647
rect 13461 23613 13495 23647
rect 14473 23613 14507 23647
rect 14657 23613 14691 23647
rect 15945 23613 15979 23647
rect 16221 23613 16255 23647
rect 16957 23613 16991 23647
rect 18613 23613 18647 23647
rect 20361 23613 20395 23647
rect 3433 23545 3467 23579
rect 4721 23545 4755 23579
rect 2145 23477 2179 23511
rect 4077 23477 4111 23511
rect 7021 23477 7055 23511
rect 19165 23477 19199 23511
rect 22109 23477 22143 23511
rect 22753 23477 22787 23511
rect 2145 23273 2179 23307
rect 3433 23273 3467 23307
rect 5641 23273 5675 23307
rect 7131 23273 7165 23307
rect 10793 23273 10827 23307
rect 16589 23273 16623 23307
rect 17877 23273 17911 23307
rect 24685 23273 24719 23307
rect 7849 23137 7883 23171
rect 11437 23137 11471 23171
rect 13645 23137 13679 23171
rect 15393 23137 15427 23171
rect 17233 23137 17267 23171
rect 19533 23137 19567 23171
rect 19809 23137 19843 23171
rect 2053 23069 2087 23103
rect 2697 23069 2731 23103
rect 7389 23069 7423 23103
rect 8401 23069 8435 23103
rect 9413 23069 9447 23103
rect 10241 23069 10275 23103
rect 10701 23069 10735 23103
rect 14381 23069 14415 23103
rect 16681 23069 16715 23103
rect 17325 23069 17359 23103
rect 17969 23069 18003 23103
rect 23765 23069 23799 23103
rect 4077 23001 4111 23035
rect 5089 23001 5123 23035
rect 8493 23001 8527 23035
rect 11529 23001 11563 23035
rect 12081 23001 12115 23035
rect 13001 23001 13035 23035
rect 13553 23001 13587 23035
rect 15117 23001 15151 23035
rect 15209 23001 15243 23035
rect 19625 23001 19659 23035
rect 2789 22933 2823 22967
rect 4629 22933 4663 22967
rect 9505 22933 9539 22967
rect 10149 22933 10183 22967
rect 14473 22933 14507 22967
rect 18797 22933 18831 22967
rect 23673 22933 23707 22967
rect 1777 22729 1811 22763
rect 3985 22729 4019 22763
rect 7113 22729 7147 22763
rect 15945 22729 15979 22763
rect 18153 22729 18187 22763
rect 7941 22661 7975 22695
rect 11805 22661 11839 22695
rect 12541 22661 12575 22695
rect 14289 22661 14323 22695
rect 14841 22661 14875 22695
rect 17049 22661 17083 22695
rect 17601 22661 17635 22695
rect 1593 22593 1627 22627
rect 2237 22593 2271 22627
rect 4905 22593 4939 22627
rect 5365 22593 5399 22627
rect 5917 22593 5951 22627
rect 7021 22593 7055 22627
rect 10517 22593 10551 22627
rect 11161 22583 11195 22617
rect 11897 22593 11931 22627
rect 13737 22593 13771 22627
rect 18245 22593 18279 22627
rect 18705 22593 18739 22627
rect 19717 22593 19751 22627
rect 28641 22593 28675 22627
rect 28733 22593 28767 22627
rect 36093 22593 36127 22627
rect 2513 22525 2547 22559
rect 7665 22525 7699 22559
rect 12449 22525 12483 22559
rect 14933 22525 14967 22559
rect 16957 22525 16991 22559
rect 29285 22525 29319 22559
rect 13001 22457 13035 22491
rect 36277 22457 36311 22491
rect 9413 22389 9447 22423
rect 10425 22389 10459 22423
rect 11069 22389 11103 22423
rect 13645 22389 13679 22423
rect 19625 22389 19659 22423
rect 20269 22389 20303 22423
rect 4248 22185 4282 22219
rect 8033 22185 8067 22219
rect 11253 22185 11287 22219
rect 12541 22185 12575 22219
rect 6285 22049 6319 22083
rect 10609 22049 10643 22083
rect 13553 22049 13587 22083
rect 13737 22049 13771 22083
rect 14473 22049 14507 22083
rect 14933 22049 14967 22083
rect 16589 22049 16623 22083
rect 1869 21981 1903 22015
rect 3985 21981 4019 22015
rect 9413 21981 9447 22015
rect 10057 21991 10091 22025
rect 10517 21981 10551 22015
rect 11161 21981 11195 22015
rect 11805 21981 11839 22015
rect 12449 21991 12483 22025
rect 13093 21981 13127 22015
rect 15485 21981 15519 22015
rect 19993 21981 20027 22015
rect 26341 21981 26375 22015
rect 6561 21913 6595 21947
rect 14841 21913 14875 21947
rect 17141 21913 17175 21947
rect 17233 21913 17267 21947
rect 18153 21913 18187 21947
rect 18245 21913 18279 21947
rect 18797 21913 18831 21947
rect 1685 21845 1719 21879
rect 2881 21845 2915 21879
rect 3341 21845 3375 21879
rect 5733 21845 5767 21879
rect 8585 21845 8619 21879
rect 9321 21845 9355 21879
rect 9965 21845 9999 21879
rect 11897 21845 11931 21879
rect 15577 21845 15611 21879
rect 20177 21845 20211 21879
rect 20729 21845 20763 21879
rect 26249 21845 26283 21879
rect 6837 21641 6871 21675
rect 10057 21641 10091 21675
rect 11989 21641 12023 21675
rect 12633 21641 12667 21675
rect 16957 21641 16991 21675
rect 7573 21573 7607 21607
rect 13737 21573 13771 21607
rect 14473 21573 14507 21607
rect 14565 21573 14599 21607
rect 15117 21573 15151 21607
rect 15577 21573 15611 21607
rect 16129 21573 16163 21607
rect 18153 21573 18187 21607
rect 1869 21505 1903 21539
rect 10149 21505 10183 21539
rect 10793 21505 10827 21539
rect 12081 21505 12115 21539
rect 12725 21505 12759 21539
rect 16865 21505 16899 21539
rect 35633 21505 35667 21539
rect 36277 21505 36311 21539
rect 3341 21437 3375 21471
rect 3617 21437 3651 21471
rect 5365 21437 5399 21471
rect 6009 21437 6043 21471
rect 7297 21437 7331 21471
rect 9321 21437 9355 21471
rect 13553 21437 13587 21471
rect 13829 21437 13863 21471
rect 16221 21437 16255 21471
rect 18705 21369 18739 21403
rect 1685 21301 1719 21335
rect 2881 21301 2915 21335
rect 10701 21301 10735 21335
rect 17601 21301 17635 21335
rect 36185 21301 36219 21335
rect 2145 21097 2179 21131
rect 10977 21097 11011 21131
rect 12265 21097 12299 21131
rect 16957 21097 16991 21131
rect 18705 21097 18739 21131
rect 9689 21029 9723 21063
rect 13461 21029 13495 21063
rect 4353 20961 4387 20995
rect 6101 20961 6135 20995
rect 10333 20961 10367 20995
rect 12909 20961 12943 20995
rect 4077 20893 4111 20927
rect 6561 20893 6595 20927
rect 9597 20893 9631 20927
rect 10425 20893 10459 20927
rect 10885 20893 10919 20927
rect 11529 20893 11563 20927
rect 12173 20893 12207 20927
rect 14473 20893 14507 20927
rect 14565 20893 14599 20927
rect 16405 20893 16439 20927
rect 16865 20893 16899 20927
rect 17509 20893 17543 20927
rect 3433 20825 3467 20859
rect 6837 20825 6871 20859
rect 8585 20825 8619 20859
rect 13001 20825 13035 20859
rect 15025 20825 15059 20859
rect 15577 20825 15611 20859
rect 15669 20825 15703 20859
rect 18061 20825 18095 20859
rect 19441 20825 19475 20859
rect 19993 20825 20027 20859
rect 20085 20825 20119 20859
rect 11621 20757 11655 20791
rect 16313 20757 16347 20791
rect 3433 20553 3467 20587
rect 10425 20553 10459 20587
rect 11069 20553 11103 20587
rect 15209 20553 15243 20587
rect 16865 20553 16899 20587
rect 20361 20553 20395 20587
rect 36001 20553 36035 20587
rect 4261 20485 4295 20519
rect 6837 20485 6871 20519
rect 12817 20485 12851 20519
rect 12909 20485 12943 20519
rect 13461 20485 13495 20519
rect 14473 20485 14507 20519
rect 1685 20417 1719 20451
rect 9321 20417 9355 20451
rect 10517 20417 10551 20451
rect 10977 20417 11011 20451
rect 12081 20417 12115 20451
rect 15301 20417 15335 20451
rect 16221 20417 16255 20451
rect 17417 20417 17451 20451
rect 20177 20417 20211 20451
rect 20821 20417 20855 20451
rect 35817 20417 35851 20451
rect 1961 20349 1995 20383
rect 5917 20349 5951 20383
rect 7297 20349 7331 20383
rect 7573 20349 7607 20383
rect 14565 20349 14599 20383
rect 19165 20349 19199 20383
rect 14013 20281 14047 20315
rect 16037 20281 16071 20315
rect 17509 20281 17543 20315
rect 9873 20213 9907 20247
rect 12173 20213 12207 20247
rect 18153 20213 18187 20247
rect 18613 20213 18647 20247
rect 35265 20213 35299 20247
rect 1685 20009 1719 20043
rect 6009 20009 6043 20043
rect 9873 20009 9907 20043
rect 14381 20009 14415 20043
rect 15117 20009 15151 20043
rect 17509 20009 17543 20043
rect 10517 19941 10551 19975
rect 12357 19941 12391 19975
rect 18797 19941 18831 19975
rect 3433 19873 3467 19907
rect 4261 19873 4295 19907
rect 4537 19873 4571 19907
rect 6745 19873 6779 19907
rect 8493 19873 8527 19907
rect 11805 19873 11839 19907
rect 12909 19873 12943 19907
rect 13553 19873 13587 19907
rect 19533 19873 19567 19907
rect 9321 19805 9355 19839
rect 9965 19805 9999 19839
rect 10609 19805 10643 19839
rect 11069 19805 11103 19839
rect 14473 19805 14507 19839
rect 15209 19805 15243 19839
rect 15853 19805 15887 19839
rect 16957 19805 16991 19839
rect 17601 19805 17635 19839
rect 18245 19805 18279 19839
rect 22477 19805 22511 19839
rect 22937 19805 22971 19839
rect 3157 19737 3191 19771
rect 7021 19737 7055 19771
rect 9229 19737 9263 19771
rect 11897 19737 11931 19771
rect 13461 19737 13495 19771
rect 19625 19737 19659 19771
rect 20177 19737 20211 19771
rect 11161 19669 11195 19703
rect 15761 19669 15795 19703
rect 16405 19669 16439 19703
rect 18153 19669 18187 19703
rect 22385 19669 22419 19703
rect 6009 19465 6043 19499
rect 11897 19465 11931 19499
rect 14933 19465 14967 19499
rect 16221 19465 16255 19499
rect 18521 19465 18555 19499
rect 3617 19397 3651 19431
rect 7757 19397 7791 19431
rect 12633 19397 12667 19431
rect 17049 19397 17083 19431
rect 19993 19397 20027 19431
rect 22201 19397 22235 19431
rect 1593 19329 1627 19363
rect 4261 19329 4295 19363
rect 6929 19329 6963 19363
rect 7021 19329 7055 19363
rect 9505 19329 9539 19363
rect 10517 19329 10551 19363
rect 10977 19329 11011 19363
rect 11805 19329 11839 19363
rect 14289 19329 14323 19363
rect 14381 19329 14415 19363
rect 15025 19329 15059 19363
rect 15669 19329 15703 19363
rect 16313 19329 16347 19363
rect 18429 19329 18463 19363
rect 19073 19329 19107 19363
rect 19165 19329 19199 19363
rect 35909 19329 35943 19363
rect 1869 19261 1903 19295
rect 4537 19261 4571 19295
rect 7481 19261 7515 19295
rect 12541 19261 12575 19295
rect 13185 19261 13219 19295
rect 16957 19261 16991 19295
rect 17233 19261 17267 19295
rect 19901 19261 19935 19295
rect 20177 19261 20211 19295
rect 21097 19261 21131 19295
rect 22109 19261 22143 19295
rect 22385 19261 22419 19295
rect 13737 19193 13771 19227
rect 10425 19125 10459 19159
rect 11069 19125 11103 19159
rect 15577 19125 15611 19159
rect 36093 19125 36127 19159
rect 1593 18921 1627 18955
rect 6837 18921 6871 18955
rect 9505 18921 9539 18955
rect 14381 18921 14415 18955
rect 16957 18921 16991 18955
rect 18245 18853 18279 18887
rect 3065 18785 3099 18819
rect 3341 18785 3375 18819
rect 5733 18785 5767 18819
rect 6009 18785 6043 18819
rect 8585 18785 8619 18819
rect 11437 18785 11471 18819
rect 13185 18785 13219 18819
rect 15485 18785 15519 18819
rect 16405 18785 16439 18819
rect 19533 18785 19567 18819
rect 21833 18785 21867 18819
rect 3985 18717 4019 18751
rect 9597 18717 9631 18751
rect 10241 18717 10275 18751
rect 10701 18717 10735 18751
rect 17417 18717 17451 18751
rect 8309 18649 8343 18683
rect 11529 18649 11563 18683
rect 12081 18649 12115 18683
rect 12541 18649 12575 18683
rect 13093 18649 13127 18683
rect 14841 18649 14875 18683
rect 15393 18649 15427 18683
rect 17601 18649 17635 18683
rect 18705 18649 18739 18683
rect 18797 18649 18831 18683
rect 19625 18649 19659 18683
rect 20545 18649 20579 18683
rect 21189 18649 21223 18683
rect 21741 18649 21775 18683
rect 10149 18581 10183 18615
rect 10793 18581 10827 18615
rect 1961 18377 1995 18411
rect 6653 18377 6687 18411
rect 18705 18377 18739 18411
rect 21281 18377 21315 18411
rect 22937 18377 22971 18411
rect 7481 18309 7515 18343
rect 12081 18309 12115 18343
rect 12633 18309 12667 18343
rect 13737 18309 13771 18343
rect 15209 18309 15243 18343
rect 15301 18309 15335 18343
rect 16957 18309 16991 18343
rect 20545 18309 20579 18343
rect 5917 18241 5951 18275
rect 6745 18241 6779 18275
rect 10333 18241 10367 18275
rect 10977 18241 11011 18275
rect 17049 18241 17083 18275
rect 19349 18241 19383 18275
rect 21373 18241 21407 18275
rect 22477 18241 22511 18275
rect 24961 18241 24995 18275
rect 25513 18241 25547 18275
rect 36093 18241 36127 18275
rect 3433 18173 3467 18207
rect 3709 18173 3743 18207
rect 5641 18173 5675 18207
rect 7205 18173 7239 18207
rect 9229 18173 9263 18207
rect 11989 18173 12023 18207
rect 13645 18173 13679 18207
rect 14657 18173 14691 18207
rect 15853 18173 15887 18207
rect 20177 18173 20211 18207
rect 20637 18173 20671 18207
rect 24869 18105 24903 18139
rect 4169 18037 4203 18071
rect 10241 18037 10275 18071
rect 11069 18037 11103 18071
rect 17877 18037 17911 18071
rect 19441 18037 19475 18071
rect 22385 18037 22419 18071
rect 36277 18037 36311 18071
rect 1856 17833 1890 17867
rect 8493 17833 8527 17867
rect 10793 17833 10827 17867
rect 16129 17833 16163 17867
rect 21925 17833 21959 17867
rect 3341 17765 3375 17799
rect 9505 17765 9539 17799
rect 17325 17765 17359 17799
rect 4445 17697 4479 17731
rect 7021 17697 7055 17731
rect 10149 17697 10183 17731
rect 11529 17697 11563 17731
rect 13369 17697 13403 17731
rect 14289 17697 14323 17731
rect 14933 17697 14967 17731
rect 20545 17697 20579 17731
rect 21189 17697 21223 17731
rect 23029 17697 23063 17731
rect 1593 17629 1627 17663
rect 6745 17629 6779 17663
rect 9597 17629 9631 17663
rect 10241 17629 10275 17663
rect 10885 17629 10919 17663
rect 16037 17629 16071 17663
rect 16681 17629 16715 17663
rect 19625 17629 19659 17663
rect 21833 17629 21867 17663
rect 4721 17561 4755 17595
rect 11621 17561 11655 17595
rect 12173 17561 12207 17595
rect 13093 17561 13127 17595
rect 13185 17561 13219 17595
rect 14841 17561 14875 17595
rect 16773 17561 16807 17595
rect 18153 17561 18187 17595
rect 21097 17561 21131 17595
rect 22569 17561 22603 17595
rect 6193 17493 6227 17527
rect 15577 17493 15611 17527
rect 18889 17493 18923 17527
rect 19533 17493 19567 17527
rect 1685 17289 1719 17323
rect 4813 17289 4847 17323
rect 6745 17289 6779 17323
rect 10333 17289 10367 17323
rect 11069 17289 11103 17323
rect 7573 17221 7607 17255
rect 11897 17221 11931 17255
rect 13093 17221 13127 17255
rect 14841 17221 14875 17255
rect 15393 17221 15427 17255
rect 20453 17221 20487 17255
rect 21005 17221 21039 17255
rect 22017 17221 22051 17255
rect 1869 17153 1903 17187
rect 2605 17153 2639 17187
rect 6009 17153 6043 17187
rect 6837 17153 6871 17187
rect 10425 17153 10459 17187
rect 10977 17153 11011 17187
rect 14381 17153 14415 17187
rect 16221 17153 16255 17187
rect 17785 17153 17819 17187
rect 18429 17153 18463 17187
rect 19073 17153 19107 17187
rect 3065 17085 3099 17119
rect 3341 17085 3375 17119
rect 7297 17085 7331 17119
rect 9321 17085 9355 17119
rect 11805 17085 11839 17119
rect 13001 17085 13035 17119
rect 13645 17085 13679 17119
rect 15485 17085 15519 17119
rect 16865 17085 16899 17119
rect 21097 17085 21131 17119
rect 2421 17017 2455 17051
rect 12357 17017 12391 17051
rect 18889 17017 18923 17051
rect 5917 16949 5951 16983
rect 14289 16949 14323 16983
rect 16129 16949 16163 16983
rect 18337 16949 18371 16983
rect 19717 16949 19751 16983
rect 3341 16745 3375 16779
rect 19533 16745 19567 16779
rect 20821 16745 20855 16779
rect 21465 16745 21499 16779
rect 7297 16677 7331 16711
rect 17417 16677 17451 16711
rect 21925 16677 21959 16711
rect 22477 16677 22511 16711
rect 1593 16609 1627 16643
rect 1869 16609 1903 16643
rect 4261 16609 4295 16643
rect 4721 16609 4755 16643
rect 9137 16609 9171 16643
rect 11437 16609 11471 16643
rect 13185 16609 13219 16643
rect 15669 16609 15703 16643
rect 15945 16609 15979 16643
rect 16865 16609 16899 16643
rect 19993 16609 20027 16643
rect 6745 16541 6779 16575
rect 7941 16541 7975 16575
rect 8493 16541 8527 16575
rect 8585 16541 8619 16575
rect 11345 16541 11379 16575
rect 12173 16541 12207 16575
rect 14841 16541 14875 16575
rect 18245 16541 18279 16575
rect 20729 16541 20763 16575
rect 4997 16473 5031 16507
rect 10885 16473 10919 16507
rect 12725 16473 12759 16507
rect 12817 16473 12851 16507
rect 15853 16473 15887 16507
rect 16957 16473 16991 16507
rect 7849 16405 7883 16439
rect 14657 16405 14691 16439
rect 18337 16405 18371 16439
rect 11897 16201 11931 16235
rect 16037 16201 16071 16235
rect 16957 16201 16991 16235
rect 22017 16201 22051 16235
rect 2881 16133 2915 16167
rect 7665 16133 7699 16167
rect 10149 16133 10183 16167
rect 12541 16133 12575 16167
rect 13277 16133 13311 16167
rect 14473 16133 14507 16167
rect 18521 16133 18555 16167
rect 19717 16133 19751 16167
rect 20361 16133 20395 16167
rect 1869 16065 1903 16099
rect 4905 16065 4939 16099
rect 5917 16065 5951 16099
rect 6009 16065 6043 16099
rect 6929 16065 6963 16099
rect 9413 16065 9447 16099
rect 10977 16065 11011 16099
rect 11805 16065 11839 16099
rect 12449 16065 12483 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 22569 16065 22603 16099
rect 26433 16065 26467 16099
rect 35725 16065 35759 16099
rect 36369 16065 36403 16099
rect 4629 15997 4663 16031
rect 6837 15997 6871 16031
rect 7389 15997 7423 16031
rect 13185 15997 13219 16031
rect 14381 15997 14415 16031
rect 15301 15997 15335 16031
rect 17969 15997 18003 16031
rect 18613 15997 18647 16031
rect 19809 15997 19843 16031
rect 26341 15997 26375 16031
rect 1685 15929 1719 15963
rect 10333 15929 10367 15963
rect 13737 15929 13771 15963
rect 19257 15929 19291 15963
rect 2329 15861 2363 15895
rect 11069 15861 11103 15895
rect 21005 15861 21039 15895
rect 36185 15861 36219 15895
rect 3341 15657 3375 15691
rect 10885 15657 10919 15691
rect 17325 15657 17359 15691
rect 18705 15657 18739 15691
rect 21649 15657 21683 15691
rect 19993 15589 20027 15623
rect 1593 15521 1627 15555
rect 8309 15521 8343 15555
rect 12541 15521 12575 15555
rect 13737 15521 13771 15555
rect 15485 15521 15519 15555
rect 20545 15521 20579 15555
rect 4261 15453 4295 15487
rect 6561 15453 6595 15487
rect 8585 15453 8619 15487
rect 9137 15453 9171 15487
rect 14749 15453 14783 15487
rect 16129 15453 16163 15487
rect 17233 15453 17267 15487
rect 18061 15453 18095 15487
rect 18613 15453 18647 15487
rect 22753 15453 22787 15487
rect 1869 15385 1903 15419
rect 4537 15385 4571 15419
rect 9413 15385 9447 15419
rect 11897 15385 11931 15419
rect 11989 15385 12023 15419
rect 13093 15385 13127 15419
rect 13185 15385 13219 15419
rect 15577 15385 15611 15419
rect 20453 15385 20487 15419
rect 22201 15385 22235 15419
rect 6009 15317 6043 15351
rect 14841 15317 14875 15351
rect 16773 15317 16807 15351
rect 17969 15317 18003 15351
rect 21097 15317 21131 15351
rect 5549 15113 5583 15147
rect 11805 15113 11839 15147
rect 18153 15113 18187 15147
rect 1593 15045 1627 15079
rect 3341 15045 3375 15079
rect 6653 15045 6687 15079
rect 10977 15045 11011 15079
rect 12817 15045 12851 15079
rect 13369 15045 13403 15079
rect 14197 15045 14231 15079
rect 15393 15045 15427 15079
rect 16957 15045 16991 15079
rect 17049 15045 17083 15079
rect 18705 15045 18739 15079
rect 19349 15045 19383 15079
rect 20085 15045 20119 15079
rect 20637 15045 20671 15079
rect 4261 14977 4295 15011
rect 6745 14977 6779 15011
rect 9965 14977 9999 15011
rect 11713 14977 11747 15011
rect 14749 14977 14783 15011
rect 18061 14977 18095 15011
rect 19257 14977 19291 15011
rect 21097 14977 21131 15011
rect 3617 14909 3651 14943
rect 7297 14909 7331 14943
rect 7573 14909 7607 14943
rect 9321 14909 9355 14943
rect 10701 14909 10735 14943
rect 11069 14909 11103 14943
rect 13461 14909 13495 14943
rect 14105 14909 14139 14943
rect 15301 14909 15335 14943
rect 15669 14909 15703 14943
rect 17233 14909 17267 14943
rect 19993 14909 20027 14943
rect 21189 14909 21223 14943
rect 22569 14909 22603 14943
rect 9873 14773 9907 14807
rect 22109 14773 22143 14807
rect 3433 14569 3467 14603
rect 4813 14569 4847 14603
rect 13001 14569 13035 14603
rect 13645 14569 13679 14603
rect 15025 14569 15059 14603
rect 16037 14569 16071 14603
rect 18797 14569 18831 14603
rect 1685 14433 1719 14467
rect 1961 14433 1995 14467
rect 8585 14433 8619 14467
rect 9137 14433 9171 14467
rect 9413 14433 9447 14467
rect 18061 14433 18095 14467
rect 19993 14433 20027 14467
rect 22385 14433 22419 14467
rect 6101 14365 6135 14399
rect 13093 14365 13127 14399
rect 13737 14365 13771 14399
rect 14473 14365 14507 14399
rect 15117 14365 15151 14399
rect 16129 14365 16163 14399
rect 36093 14365 36127 14399
rect 6561 14297 6595 14331
rect 8309 14297 8343 14331
rect 11437 14297 11471 14331
rect 11989 14297 12023 14331
rect 12081 14297 12115 14331
rect 17141 14297 17175 14331
rect 17693 14297 17727 14331
rect 17785 14297 17819 14331
rect 20085 14297 20119 14331
rect 20637 14297 20671 14331
rect 21097 14297 21131 14331
rect 21649 14297 21683 14331
rect 21741 14297 21775 14331
rect 22477 14297 22511 14331
rect 23029 14297 23063 14331
rect 10885 14229 10919 14263
rect 35541 14229 35575 14263
rect 36277 14229 36311 14263
rect 11069 14025 11103 14059
rect 12081 14025 12115 14059
rect 21097 14025 21131 14059
rect 1961 13957 1995 13991
rect 7389 13957 7423 13991
rect 9873 13957 9907 13991
rect 12817 13957 12851 13991
rect 14289 13957 14323 13991
rect 14841 13957 14875 13991
rect 15485 13957 15519 13991
rect 16957 13957 16991 13991
rect 17049 13957 17083 13991
rect 18521 13957 18555 13991
rect 20361 13957 20395 13991
rect 22109 13957 22143 13991
rect 22201 13957 22235 13991
rect 23305 13957 23339 13991
rect 1685 13889 1719 13923
rect 4261 13889 4295 13923
rect 9965 13889 9999 13923
rect 10977 13889 11011 13923
rect 11989 13889 12023 13923
rect 18613 13889 18647 13923
rect 19257 13889 19291 13923
rect 21005 13889 21039 13923
rect 22753 13889 22787 13923
rect 23397 13889 23431 13923
rect 23857 13889 23891 13923
rect 3433 13821 3467 13855
rect 4537 13821 4571 13855
rect 6009 13821 6043 13855
rect 7113 13821 7147 13855
rect 9137 13821 9171 13855
rect 12725 13821 12759 13855
rect 13369 13821 13403 13855
rect 14197 13821 14231 13855
rect 15393 13821 15427 13855
rect 16037 13821 16071 13855
rect 17601 13821 17635 13855
rect 19809 13821 19843 13855
rect 20453 13821 20487 13855
rect 6653 13753 6687 13787
rect 10517 13685 10551 13719
rect 19165 13685 19199 13719
rect 1685 13481 1719 13515
rect 9781 13481 9815 13515
rect 13645 13481 13679 13515
rect 15209 13481 15243 13515
rect 16221 13481 16255 13515
rect 18061 13481 18095 13515
rect 19441 13481 19475 13515
rect 20177 13481 20211 13515
rect 21833 13481 21867 13515
rect 22477 13481 22511 13515
rect 5641 13413 5675 13447
rect 10425 13413 10459 13447
rect 14565 13413 14599 13447
rect 20821 13413 20855 13447
rect 3433 13345 3467 13379
rect 6561 13345 6595 13379
rect 8585 13345 8619 13379
rect 4353 13277 4387 13311
rect 9873 13277 9907 13311
rect 10517 13277 10551 13311
rect 11437 13277 11471 13311
rect 13553 13277 13587 13311
rect 14473 13277 14507 13311
rect 15117 13277 15151 13311
rect 16313 13277 16347 13311
rect 17969 13277 18003 13311
rect 18797 13277 18831 13311
rect 20085 13277 20119 13311
rect 21925 13277 21959 13311
rect 22569 13277 22603 13311
rect 23029 13277 23063 13311
rect 35909 13277 35943 13311
rect 3157 13209 3191 13243
rect 6837 13209 6871 13243
rect 9137 13209 9171 13243
rect 12173 13209 12207 13243
rect 12265 13209 12299 13243
rect 12817 13209 12851 13243
rect 16773 13209 16807 13243
rect 17325 13209 17359 13243
rect 17417 13209 17451 13243
rect 18705 13209 18739 13243
rect 11529 13141 11563 13175
rect 36093 13141 36127 13175
rect 5825 12937 5859 12971
rect 9965 12937 9999 12971
rect 10609 12937 10643 12971
rect 12449 12937 12483 12971
rect 20821 12937 20855 12971
rect 22109 12937 22143 12971
rect 4353 12869 4387 12903
rect 9321 12869 9355 12903
rect 13185 12869 13219 12903
rect 14381 12869 14415 12903
rect 16129 12869 16163 12903
rect 17049 12869 17083 12903
rect 19441 12869 19475 12903
rect 19533 12869 19567 12903
rect 3617 12801 3651 12835
rect 4077 12801 4111 12835
rect 6837 12801 6871 12835
rect 10057 12801 10091 12835
rect 10517 12801 10551 12835
rect 11713 12801 11747 12835
rect 12357 12801 12391 12835
rect 18061 12801 18095 12835
rect 20085 12801 20119 12835
rect 20913 12801 20947 12835
rect 35633 12801 35667 12835
rect 36277 12801 36311 12835
rect 1593 12733 1627 12767
rect 3341 12733 3375 12767
rect 7297 12733 7331 12767
rect 7573 12733 7607 12767
rect 13093 12733 13127 12767
rect 14289 12733 14323 12767
rect 14565 12733 14599 12767
rect 15945 12733 15979 12767
rect 16221 12733 16255 12767
rect 16957 12733 16991 12767
rect 17233 12733 17267 12767
rect 19257 12733 19291 12767
rect 6653 12665 6687 12699
rect 11805 12665 11839 12699
rect 13645 12665 13679 12699
rect 21465 12665 21499 12699
rect 36093 12665 36127 12699
rect 20177 12597 20211 12631
rect 1685 12393 1719 12427
rect 9321 12393 9355 12427
rect 9965 12393 9999 12427
rect 10609 12393 10643 12427
rect 13645 12393 13679 12427
rect 14381 12393 14415 12427
rect 16681 12393 16715 12427
rect 18521 12393 18555 12427
rect 3157 12257 3191 12291
rect 6009 12257 6043 12291
rect 8585 12257 8619 12291
rect 11529 12257 11563 12291
rect 11805 12257 11839 12291
rect 14933 12257 14967 12291
rect 15577 12257 15611 12291
rect 17233 12257 17267 12291
rect 17877 12257 17911 12291
rect 3433 12189 3467 12223
rect 9413 12189 9447 12223
rect 10057 12189 10091 12223
rect 10517 12189 10551 12223
rect 14473 12189 14507 12223
rect 16773 12189 16807 12223
rect 5733 12121 5767 12155
rect 6561 12121 6595 12155
rect 8309 12121 8343 12155
rect 11713 12121 11747 12155
rect 12449 12121 12483 12155
rect 13001 12121 13035 12155
rect 13093 12121 13127 12155
rect 15485 12121 15519 12155
rect 17792 12121 17826 12155
rect 19533 12121 19567 12155
rect 20085 12121 20119 12155
rect 20177 12121 20211 12155
rect 20729 12121 20763 12155
rect 4261 12053 4295 12087
rect 1593 11849 1627 11883
rect 6745 11849 6779 11883
rect 10057 11849 10091 11883
rect 12725 11849 12759 11883
rect 14933 11849 14967 11883
rect 15577 11849 15611 11883
rect 19717 11849 19751 11883
rect 20361 11849 20395 11883
rect 7757 11781 7791 11815
rect 10885 11781 10919 11815
rect 17325 11781 17359 11815
rect 17417 11781 17451 11815
rect 6653 11713 6687 11747
rect 10241 11713 10275 11747
rect 11161 11713 11195 11747
rect 11713 11713 11747 11747
rect 12633 11713 12667 11747
rect 13277 11713 13311 11747
rect 14197 11713 14231 11747
rect 14841 11713 14875 11747
rect 15485 11713 15519 11747
rect 16221 11713 16255 11747
rect 16313 11713 16347 11747
rect 18613 11713 18647 11747
rect 19073 11713 19107 11747
rect 19809 11713 19843 11747
rect 3065 11645 3099 11679
rect 3341 11645 3375 11679
rect 3985 11645 4019 11679
rect 4261 11645 4295 11679
rect 6009 11645 6043 11679
rect 7481 11645 7515 11679
rect 9505 11645 9539 11679
rect 11897 11645 11931 11679
rect 13369 11577 13403 11611
rect 17877 11577 17911 11611
rect 14289 11509 14323 11543
rect 18521 11509 18555 11543
rect 3433 11305 3467 11339
rect 4261 11305 4295 11339
rect 10885 11305 10919 11339
rect 12725 11305 12759 11339
rect 13369 11305 13403 11339
rect 19441 11305 19475 11339
rect 36277 11237 36311 11271
rect 6009 11169 6043 11203
rect 8585 11169 8619 11203
rect 9137 11169 9171 11203
rect 14841 11169 14875 11203
rect 15853 11169 15887 11203
rect 16773 11169 16807 11203
rect 17417 11169 17451 11203
rect 1685 11101 1719 11135
rect 6561 11101 6595 11135
rect 11897 11101 11931 11135
rect 12633 11101 12667 11135
rect 13277 11101 13311 11135
rect 36093 11101 36127 11135
rect 1961 11033 1995 11067
rect 5733 11033 5767 11067
rect 8309 11033 8343 11067
rect 9413 11033 9447 11067
rect 11621 11033 11655 11067
rect 14381 11033 14415 11067
rect 14473 11033 14507 11067
rect 16037 11033 16071 11067
rect 16129 11033 16163 11067
rect 16865 11033 16899 11067
rect 17969 11033 18003 11067
rect 18061 11033 18095 11067
rect 18613 11033 18647 11067
rect 3893 10761 3927 10795
rect 6929 10761 6963 10795
rect 10149 10761 10183 10795
rect 19625 10761 19659 10795
rect 12265 10693 12299 10727
rect 14749 10693 14783 10727
rect 14841 10693 14875 10727
rect 16037 10693 16071 10727
rect 17049 10693 17083 10727
rect 2605 10625 2639 10659
rect 4997 10625 5031 10659
rect 6837 10625 6871 10659
rect 7573 10625 7607 10659
rect 10241 10625 10275 10659
rect 10885 10625 10919 10659
rect 13093 10625 13127 10659
rect 13737 10625 13771 10659
rect 17601 10625 17635 10659
rect 18889 10625 18923 10659
rect 2145 10557 2179 10591
rect 7849 10557 7883 10591
rect 9597 10557 9631 10591
rect 11713 10557 11747 10591
rect 12357 10557 12391 10591
rect 15669 10557 15703 10591
rect 16129 10557 16163 10591
rect 16957 10557 16991 10591
rect 14289 10489 14323 10523
rect 4905 10421 4939 10455
rect 6009 10421 6043 10455
rect 10793 10421 10827 10455
rect 13001 10421 13035 10455
rect 13645 10421 13679 10455
rect 19073 10421 19107 10455
rect 4813 10217 4847 10251
rect 8493 10217 8527 10251
rect 15853 10217 15887 10251
rect 4077 10149 4111 10183
rect 12725 10149 12759 10183
rect 1593 10081 1627 10115
rect 1869 10081 1903 10115
rect 3341 10081 3375 10115
rect 5733 10081 5767 10115
rect 9321 10081 9355 10115
rect 11805 10081 11839 10115
rect 12081 10081 12115 10115
rect 13277 10081 13311 10115
rect 14933 10081 14967 10115
rect 4261 10013 4295 10047
rect 4997 10013 5031 10047
rect 8401 10013 8435 10047
rect 9413 10013 9447 10047
rect 10425 10013 10459 10047
rect 15761 10013 15795 10047
rect 6009 9945 6043 9979
rect 10149 9945 10183 9979
rect 11989 9945 12023 9979
rect 13185 9945 13219 9979
rect 14289 9945 14323 9979
rect 14841 9945 14875 9979
rect 7481 9877 7515 9911
rect 10885 9877 10919 9911
rect 16497 9877 16531 9911
rect 17049 9877 17083 9911
rect 8309 9673 8343 9707
rect 3065 9605 3099 9639
rect 9413 9605 9447 9639
rect 12909 9605 12943 9639
rect 14841 9605 14875 9639
rect 6561 9537 6595 9571
rect 9321 9537 9355 9571
rect 10241 9537 10275 9571
rect 12173 9537 12207 9571
rect 13001 9537 13035 9571
rect 13921 9537 13955 9571
rect 14933 9537 14967 9571
rect 1593 9469 1627 9503
rect 3341 9469 3375 9503
rect 4261 9469 4295 9503
rect 4537 9469 4571 9503
rect 6837 9469 6871 9503
rect 10425 9469 10459 9503
rect 12265 9469 12299 9503
rect 6009 9333 6043 9367
rect 8769 9333 8803 9367
rect 13829 9333 13863 9367
rect 15853 9333 15887 9367
rect 3433 9129 3467 9163
rect 6561 9129 6595 9163
rect 7757 9129 7791 9163
rect 8493 9129 8527 9163
rect 10241 9129 10275 9163
rect 13277 9129 13311 9163
rect 14933 9129 14967 9163
rect 9597 9061 9631 9095
rect 10885 9061 10919 9095
rect 14289 9061 14323 9095
rect 36093 9061 36127 9095
rect 1685 8993 1719 9027
rect 4261 8993 4295 9027
rect 6009 8993 6043 9027
rect 12633 8993 12667 9027
rect 6653 8925 6687 8959
rect 7297 8925 7331 8959
rect 7941 8925 7975 8959
rect 8585 8925 8619 8959
rect 9689 8925 9723 8959
rect 10149 8925 10183 8959
rect 10977 8925 11011 8959
rect 11897 8925 11931 8959
rect 12541 8925 12575 8959
rect 13185 8925 13219 8959
rect 1961 8857 1995 8891
rect 5733 8857 5767 8891
rect 11989 8857 12023 8891
rect 35633 8857 35667 8891
rect 36277 8857 36311 8891
rect 7205 8789 7239 8823
rect 15393 8789 15427 8823
rect 2053 8585 2087 8619
rect 5733 8585 5767 8619
rect 7757 8585 7791 8619
rect 9321 8585 9355 8619
rect 11161 8585 11195 8619
rect 11805 8585 11839 8619
rect 12817 8585 12851 8619
rect 13461 8585 13495 8619
rect 14013 8585 14047 8619
rect 14565 8585 14599 8619
rect 16957 8585 16991 8619
rect 2605 8517 2639 8551
rect 4353 8517 4387 8551
rect 8401 8517 8435 8551
rect 10425 8517 10459 8551
rect 10517 8517 10551 8551
rect 2145 8449 2179 8483
rect 4997 8449 5031 8483
rect 5641 8449 5675 8483
rect 7205 8449 7239 8483
rect 7849 8449 7883 8483
rect 8493 8449 8527 8483
rect 9413 8449 9447 8483
rect 11713 8449 11747 8483
rect 17049 8449 17083 8483
rect 9873 8381 9907 8415
rect 4813 8313 4847 8347
rect 7113 8245 7147 8279
rect 3433 8041 3467 8075
rect 5733 8041 5767 8075
rect 10885 8041 10919 8075
rect 11529 8041 11563 8075
rect 13461 8041 13495 8075
rect 36185 8041 36219 8075
rect 7481 7973 7515 8007
rect 1685 7905 1719 7939
rect 1961 7905 1995 7939
rect 4261 7905 4295 7939
rect 12817 7905 12851 7939
rect 3985 7837 4019 7871
rect 7021 7837 7055 7871
rect 8585 7837 8619 7871
rect 9413 7837 9447 7871
rect 10793 7837 10827 7871
rect 11437 7837 11471 7871
rect 9689 7769 9723 7803
rect 35633 7769 35667 7803
rect 36277 7769 36311 7803
rect 8493 7701 8527 7735
rect 12173 7701 12207 7735
rect 3801 7497 3835 7531
rect 6653 7497 6687 7531
rect 7849 7497 7883 7531
rect 8401 7497 8435 7531
rect 12449 7497 12483 7531
rect 3341 7361 3375 7395
rect 5549 7361 5583 7395
rect 6561 7361 6595 7395
rect 8309 7361 8343 7395
rect 9229 7361 9263 7395
rect 11989 7361 12023 7395
rect 3065 7293 3099 7327
rect 5273 7293 5307 7327
rect 9413 7293 9447 7327
rect 1593 7225 1627 7259
rect 7297 7225 7331 7259
rect 10609 7225 10643 7259
rect 11805 7157 11839 7191
rect 1948 6953 1982 6987
rect 1685 6817 1719 6851
rect 4077 6817 4111 6851
rect 5273 6817 5307 6851
rect 5917 6817 5951 6851
rect 7481 6817 7515 6851
rect 8585 6817 8619 6851
rect 10333 6817 10367 6851
rect 11069 6817 11103 6851
rect 4721 6749 4755 6783
rect 5365 6749 5399 6783
rect 6009 6749 6043 6783
rect 9137 6749 9171 6783
rect 22385 6749 22419 6783
rect 4629 6681 4663 6715
rect 12633 6681 12667 6715
rect 13185 6681 13219 6715
rect 13277 6681 13311 6715
rect 3433 6613 3467 6647
rect 7021 6613 7055 6647
rect 9689 6613 9723 6647
rect 22477 6613 22511 6647
rect 1685 6409 1719 6443
rect 4261 6409 4295 6443
rect 5917 6409 5951 6443
rect 6561 6409 6595 6443
rect 7481 6409 7515 6443
rect 8033 6409 8067 6443
rect 9045 6409 9079 6443
rect 9597 6409 9631 6443
rect 13001 6409 13035 6443
rect 3157 6341 3191 6375
rect 4905 6341 4939 6375
rect 10057 6341 10091 6375
rect 3433 6273 3467 6307
rect 4169 6273 4203 6307
rect 4813 6273 4847 6307
rect 22109 6273 22143 6307
rect 22753 6273 22787 6307
rect 22293 6137 22327 6171
rect 1685 5865 1719 5899
rect 2973 5865 3007 5899
rect 4077 5865 4111 5899
rect 5181 5865 5215 5899
rect 6101 5865 6135 5899
rect 7849 5865 7883 5899
rect 6653 5797 6687 5831
rect 7297 5797 7331 5831
rect 1777 5661 1811 5695
rect 2421 5661 2455 5695
rect 3065 5661 3099 5695
rect 3985 5661 4019 5695
rect 36093 5661 36127 5695
rect 2329 5593 2363 5627
rect 4629 5593 4663 5627
rect 35541 5593 35575 5627
rect 36277 5525 36311 5559
rect 2697 5321 2731 5355
rect 4629 5321 4663 5355
rect 5181 5321 5215 5355
rect 5733 5321 5767 5355
rect 17693 5321 17727 5355
rect 1869 5185 1903 5219
rect 2605 5185 2639 5219
rect 3249 5185 3283 5219
rect 4077 5185 4111 5219
rect 16957 5185 16991 5219
rect 3341 5049 3375 5083
rect 1685 4981 1719 5015
rect 3893 4981 3927 5015
rect 17141 4981 17175 5015
rect 2053 4777 2087 4811
rect 2697 4777 2731 4811
rect 3341 4777 3375 4811
rect 3985 4777 4019 4811
rect 4721 4777 4755 4811
rect 5273 4777 5307 4811
rect 1961 4573 1995 4607
rect 2789 4573 2823 4607
rect 9321 4573 9355 4607
rect 36093 4573 36127 4607
rect 9229 4437 9263 4471
rect 36277 4437 36311 4471
rect 2605 4233 2639 4267
rect 3157 4233 3191 4267
rect 1961 4097 1995 4131
rect 2421 4097 2455 4131
rect 3893 4097 3927 4131
rect 25881 4097 25915 4131
rect 26525 4097 26559 4131
rect 1869 4029 1903 4063
rect 26065 3961 26099 3995
rect 2421 3689 2455 3723
rect 1869 3485 1903 3519
rect 19441 3485 19475 3519
rect 35633 3485 35667 3519
rect 36277 3485 36311 3519
rect 36093 3417 36127 3451
rect 1685 3349 1719 3383
rect 19533 3349 19567 3383
rect 35449 3145 35483 3179
rect 36185 3145 36219 3179
rect 1869 3009 1903 3043
rect 7297 3009 7331 3043
rect 18613 3009 18647 3043
rect 34897 3009 34931 3043
rect 35541 3009 35575 3043
rect 36277 3009 36311 3043
rect 2421 2873 2455 2907
rect 1685 2805 1719 2839
rect 7481 2805 7515 2839
rect 18797 2805 18831 2839
rect 27169 2805 27203 2839
rect 30389 2805 30423 2839
rect 4215 2601 4249 2635
rect 13001 2601 13035 2635
rect 14473 2601 14507 2635
rect 29837 2601 29871 2635
rect 30573 2601 30607 2635
rect 32413 2601 32447 2635
rect 34989 2601 35023 2635
rect 2421 2533 2455 2567
rect 11989 2533 12023 2567
rect 16313 2533 16347 2567
rect 27169 2533 27203 2567
rect 33885 2533 33919 2567
rect 1869 2397 1903 2431
rect 2605 2397 2639 2431
rect 3985 2397 4019 2431
rect 5549 2397 5583 2431
rect 6837 2397 6871 2431
rect 7389 2397 7423 2431
rect 7849 2397 7883 2431
rect 10057 2397 10091 2431
rect 13185 2397 13219 2431
rect 13645 2397 13679 2431
rect 14289 2397 14323 2431
rect 14933 2397 14967 2431
rect 17509 2397 17543 2431
rect 19441 2397 19475 2431
rect 20729 2397 20763 2431
rect 22661 2397 22695 2431
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 30665 2397 30699 2431
rect 35541 2397 35575 2431
rect 9321 2329 9355 2363
rect 9873 2329 9907 2363
rect 11805 2329 11839 2363
rect 16129 2329 16163 2363
rect 16865 2329 16899 2363
rect 27353 2329 27387 2363
rect 29929 2329 29963 2363
rect 31769 2329 31803 2363
rect 32505 2329 32539 2363
rect 33149 2329 33183 2363
rect 33701 2329 33735 2363
rect 1685 2261 1719 2295
rect 3341 2261 3375 2295
rect 5365 2261 5399 2295
rect 6653 2261 6687 2295
rect 8033 2261 8067 2295
rect 11069 2261 11103 2295
rect 17693 2261 17727 2295
rect 19625 2261 19659 2295
rect 20913 2261 20947 2295
rect 22845 2261 22879 2295
rect 24777 2261 24811 2295
rect 26065 2261 26099 2295
rect 29101 2261 29135 2295
rect 35725 2261 35759 2295
rect 36369 2261 36403 2295
<< metal1 >>
rect 1104 37562 36892 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 36892 37562
rect 1104 37488 36892 37510
rect 14461 37451 14519 37457
rect 14461 37417 14473 37451
rect 14507 37448 14519 37451
rect 14826 37448 14832 37460
rect 14507 37420 14832 37448
rect 14507 37417 14519 37420
rect 14461 37411 14519 37417
rect 14826 37408 14832 37420
rect 14884 37408 14890 37460
rect 26418 37408 26424 37460
rect 26476 37448 26482 37460
rect 26513 37451 26571 37457
rect 26513 37448 26525 37451
rect 26476 37420 26525 37448
rect 26476 37408 26482 37420
rect 26513 37417 26525 37420
rect 26559 37417 26571 37451
rect 26513 37411 26571 37417
rect 32493 37451 32551 37457
rect 32493 37417 32505 37451
rect 32539 37448 32551 37451
rect 32858 37448 32864 37460
rect 32539 37420 32864 37448
rect 32539 37417 32551 37420
rect 32493 37411 32551 37417
rect 5905 37315 5963 37321
rect 5905 37312 5917 37315
rect 5460 37284 5917 37312
rect 2314 37244 2320 37256
rect 2275 37216 2320 37244
rect 2314 37204 2320 37216
rect 2372 37204 2378 37256
rect 3053 37247 3111 37253
rect 3053 37213 3065 37247
rect 3099 37244 3111 37247
rect 3234 37244 3240 37256
rect 3099 37216 3240 37244
rect 3099 37213 3111 37216
rect 3053 37207 3111 37213
rect 3234 37204 3240 37216
rect 3292 37204 3298 37256
rect 4246 37244 4252 37256
rect 4207 37216 4252 37244
rect 4246 37204 4252 37216
rect 4304 37204 4310 37256
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5460 37253 5488 37284
rect 5905 37281 5917 37284
rect 5951 37281 5963 37315
rect 5905 37275 5963 37281
rect 6733 37315 6791 37321
rect 6733 37281 6745 37315
rect 6779 37312 6791 37315
rect 7098 37312 7104 37324
rect 6779 37284 7104 37312
rect 6779 37281 6791 37284
rect 6733 37275 6791 37281
rect 7098 37272 7104 37284
rect 7156 37312 7162 37324
rect 7469 37315 7527 37321
rect 7156 37284 7328 37312
rect 7156 37272 7162 37284
rect 7300 37253 7328 37284
rect 7469 37281 7481 37315
rect 7515 37312 7527 37315
rect 16114 37312 16120 37324
rect 7515 37284 16120 37312
rect 7515 37281 7527 37284
rect 7469 37275 7527 37281
rect 16114 37272 16120 37284
rect 16172 37312 16178 37324
rect 26418 37312 26424 37324
rect 16172 37284 26424 37312
rect 16172 37272 16178 37284
rect 26418 37272 26424 37284
rect 26476 37272 26482 37324
rect 26528 37312 26556 37411
rect 32858 37408 32864 37420
rect 32916 37408 32922 37460
rect 34146 37408 34152 37460
rect 34204 37448 34210 37460
rect 34241 37451 34299 37457
rect 34241 37448 34253 37451
rect 34204 37420 34253 37448
rect 34204 37408 34210 37420
rect 34241 37417 34253 37420
rect 34287 37417 34299 37451
rect 34241 37411 34299 37417
rect 32876 37380 32904 37408
rect 32876 37352 33088 37380
rect 27157 37315 27215 37321
rect 27157 37312 27169 37315
rect 26528 37284 27169 37312
rect 27157 37281 27169 37284
rect 27203 37281 27215 37315
rect 32950 37312 32956 37324
rect 32911 37284 32956 37312
rect 27157 37275 27215 37281
rect 32950 37272 32956 37284
rect 33008 37272 33014 37324
rect 33060 37312 33088 37352
rect 34256 37312 34284 37411
rect 33060 37284 33180 37312
rect 34256 37284 34560 37312
rect 5445 37247 5503 37253
rect 5445 37244 5457 37247
rect 5224 37216 5457 37244
rect 5224 37204 5230 37216
rect 5445 37213 5457 37216
rect 5491 37213 5503 37247
rect 5445 37207 5503 37213
rect 7285 37247 7343 37253
rect 7285 37213 7297 37247
rect 7331 37213 7343 37247
rect 9398 37244 9404 37256
rect 9359 37216 9404 37244
rect 7285 37207 7343 37213
rect 9398 37204 9404 37216
rect 9456 37204 9462 37256
rect 10686 37244 10692 37256
rect 10647 37216 10692 37244
rect 10686 37204 10692 37216
rect 10744 37204 10750 37256
rect 10778 37204 10784 37256
rect 10836 37244 10842 37256
rect 11701 37247 11759 37253
rect 11701 37244 11713 37247
rect 10836 37216 11713 37244
rect 10836 37204 10842 37216
rect 11701 37213 11713 37216
rect 11747 37213 11759 37247
rect 11701 37207 11759 37213
rect 13725 37247 13783 37253
rect 13725 37213 13737 37247
rect 13771 37244 13783 37247
rect 13998 37244 14004 37256
rect 13771 37216 14004 37244
rect 13771 37213 13783 37216
rect 13725 37207 13783 37213
rect 13998 37204 14004 37216
rect 14056 37204 14062 37256
rect 14826 37204 14832 37256
rect 14884 37244 14890 37256
rect 15105 37247 15163 37253
rect 15105 37244 15117 37247
rect 14884 37216 15117 37244
rect 14884 37204 14890 37216
rect 15105 37213 15117 37216
rect 15151 37213 15163 37247
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 15105 37207 15163 37213
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37244 18383 37247
rect 18785 37247 18843 37253
rect 18785 37244 18797 37247
rect 18371 37216 18797 37244
rect 18371 37213 18383 37216
rect 18325 37207 18383 37213
rect 18785 37213 18797 37216
rect 18831 37213 18843 37247
rect 18785 37207 18843 37213
rect 18874 37204 18880 37256
rect 18932 37244 18938 37256
rect 20073 37247 20131 37253
rect 20073 37244 20085 37247
rect 18932 37216 20085 37244
rect 18932 37204 18938 37216
rect 20073 37213 20085 37216
rect 20119 37213 20131 37247
rect 22002 37244 22008 37256
rect 21963 37216 22008 37244
rect 20073 37207 20131 37213
rect 22002 37204 22008 37216
rect 22060 37204 22066 37256
rect 22833 37247 22891 37253
rect 22833 37213 22845 37247
rect 22879 37244 22891 37247
rect 23290 37244 23296 37256
rect 22879 37216 23296 37244
rect 22879 37213 22891 37216
rect 22833 37207 22891 37213
rect 23290 37204 23296 37216
rect 23348 37204 23354 37256
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 27430 37244 27436 37256
rect 27391 37216 27436 37244
rect 27430 37204 27436 37216
rect 27488 37204 27494 37256
rect 28442 37244 28448 37256
rect 28403 37216 28448 37244
rect 28442 37204 28448 37216
rect 28500 37204 28506 37256
rect 29086 37204 29092 37256
rect 29144 37244 29150 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 29144 37216 29745 37244
rect 29144 37204 29150 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 31018 37244 31024 37256
rect 30979 37216 31024 37244
rect 29733 37207 29791 37213
rect 31018 37204 31024 37216
rect 31076 37204 31082 37256
rect 33152 37253 33180 37284
rect 33137 37247 33195 37253
rect 33137 37213 33149 37247
rect 33183 37213 33195 37247
rect 34532 37244 34560 37284
rect 34790 37272 34796 37324
rect 34848 37312 34854 37324
rect 34885 37315 34943 37321
rect 34885 37312 34897 37315
rect 34848 37284 34897 37312
rect 34848 37272 34854 37284
rect 34885 37281 34897 37284
rect 34931 37281 34943 37315
rect 34885 37275 34943 37281
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34532 37216 35081 37244
rect 33137 37207 33195 37213
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 35618 37204 35624 37256
rect 35676 37244 35682 37256
rect 36081 37247 36139 37253
rect 36081 37244 36093 37247
rect 35676 37216 36093 37244
rect 35676 37204 35682 37216
rect 36081 37213 36093 37216
rect 36127 37213 36139 37247
rect 36081 37207 36139 37213
rect 2958 37136 2964 37188
rect 3016 37176 3022 37188
rect 3016 37148 5304 37176
rect 3016 37136 3022 37148
rect 1946 37068 1952 37120
rect 2004 37108 2010 37120
rect 2133 37111 2191 37117
rect 2133 37108 2145 37111
rect 2004 37080 2145 37108
rect 2004 37068 2010 37080
rect 2133 37077 2145 37080
rect 2179 37077 2191 37111
rect 2866 37108 2872 37120
rect 2827 37080 2872 37108
rect 2133 37071 2191 37077
rect 2866 37068 2872 37080
rect 2924 37068 2930 37120
rect 3878 37068 3884 37120
rect 3936 37108 3942 37120
rect 5276 37117 5304 37148
rect 4065 37111 4123 37117
rect 4065 37108 4077 37111
rect 3936 37080 4077 37108
rect 3936 37068 3942 37080
rect 4065 37077 4077 37080
rect 4111 37077 4123 37111
rect 4065 37071 4123 37077
rect 5261 37111 5319 37117
rect 5261 37077 5273 37111
rect 5307 37077 5319 37111
rect 5261 37071 5319 37077
rect 8386 37068 8392 37120
rect 8444 37108 8450 37120
rect 9217 37111 9275 37117
rect 9217 37108 9229 37111
rect 8444 37080 9229 37108
rect 8444 37068 8450 37080
rect 9217 37077 9229 37080
rect 9263 37077 9275 37111
rect 9217 37071 9275 37077
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10505 37111 10563 37117
rect 10505 37108 10517 37111
rect 10376 37080 10517 37108
rect 10376 37068 10382 37080
rect 10505 37077 10517 37080
rect 10551 37077 10563 37111
rect 10505 37071 10563 37077
rect 11606 37068 11612 37120
rect 11664 37108 11670 37120
rect 11885 37111 11943 37117
rect 11885 37108 11897 37111
rect 11664 37080 11897 37108
rect 11664 37068 11670 37080
rect 11885 37077 11897 37080
rect 11931 37077 11943 37111
rect 13538 37108 13544 37120
rect 13499 37080 13544 37108
rect 11885 37071 11943 37077
rect 13538 37068 13544 37080
rect 13596 37068 13602 37120
rect 15010 37108 15016 37120
rect 14971 37080 15016 37108
rect 15010 37068 15016 37080
rect 15068 37068 15074 37120
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16816 37080 17049 37108
rect 16816 37068 16822 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 18138 37108 18144 37120
rect 18099 37080 18144 37108
rect 17037 37071 17095 37077
rect 18138 37068 18144 37080
rect 18196 37068 18202 37120
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 21266 37068 21272 37120
rect 21324 37108 21330 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 21324 37080 22201 37108
rect 21324 37068 21330 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 23198 37068 23204 37120
rect 23256 37108 23262 37120
rect 23477 37111 23535 37117
rect 23477 37108 23489 37111
rect 23256 37080 23489 37108
rect 23256 37068 23262 37080
rect 23477 37077 23489 37080
rect 23523 37077 23535 37111
rect 23477 37071 23535 37077
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24544 37080 24777 37108
rect 24544 37068 24550 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 28629 37111 28687 37117
rect 28629 37108 28641 37111
rect 27764 37080 28641 37108
rect 27764 37068 27770 37080
rect 28629 37077 28641 37080
rect 28675 37077 28687 37111
rect 28629 37071 28687 37077
rect 29638 37068 29644 37120
rect 29696 37108 29702 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29696 37080 29929 37108
rect 29696 37068 29702 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 30926 37068 30932 37120
rect 30984 37108 30990 37120
rect 31205 37111 31263 37117
rect 31205 37108 31217 37111
rect 30984 37080 31217 37108
rect 30984 37068 30990 37080
rect 31205 37077 31217 37080
rect 31251 37077 31263 37111
rect 31205 37071 31263 37077
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36265 37111 36323 37117
rect 36265 37108 36277 37111
rect 36136 37080 36277 37108
rect 36136 37068 36142 37080
rect 36265 37077 36277 37080
rect 36311 37077 36323 37111
rect 36265 37071 36323 37077
rect 1104 37018 36892 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 36892 37018
rect 1104 36944 36892 36966
rect 4246 36864 4252 36916
rect 4304 36904 4310 36916
rect 4304 36876 6914 36904
rect 4304 36864 4310 36876
rect 1670 36836 1676 36848
rect 1631 36808 1676 36836
rect 1670 36796 1676 36808
rect 1728 36836 1734 36848
rect 2317 36839 2375 36845
rect 2317 36836 2329 36839
rect 1728 36808 2329 36836
rect 1728 36796 1734 36808
rect 2317 36805 2329 36808
rect 2363 36805 2375 36839
rect 6886 36836 6914 36876
rect 10686 36864 10692 36916
rect 10744 36904 10750 36916
rect 11701 36907 11759 36913
rect 11701 36904 11713 36907
rect 10744 36876 11713 36904
rect 10744 36864 10750 36876
rect 11701 36873 11713 36876
rect 11747 36873 11759 36907
rect 11701 36867 11759 36873
rect 27341 36907 27399 36913
rect 27341 36873 27353 36907
rect 27387 36904 27399 36907
rect 28442 36904 28448 36916
rect 27387 36876 28448 36904
rect 27387 36873 27399 36876
rect 27341 36867 27399 36873
rect 28442 36864 28448 36876
rect 28500 36864 28506 36916
rect 29086 36904 29092 36916
rect 29047 36876 29092 36904
rect 29086 36864 29092 36876
rect 29144 36864 29150 36916
rect 31297 36907 31355 36913
rect 31297 36873 31309 36907
rect 31343 36873 31355 36907
rect 35526 36904 35532 36916
rect 35487 36876 35532 36904
rect 31297 36867 31355 36873
rect 12250 36836 12256 36848
rect 6886 36808 12256 36836
rect 2317 36799 2375 36805
rect 12250 36796 12256 36808
rect 12308 36796 12314 36848
rect 27430 36796 27436 36848
rect 27488 36836 27494 36848
rect 27488 36808 31156 36836
rect 27488 36796 27494 36808
rect 10870 36728 10876 36780
rect 10928 36768 10934 36780
rect 11885 36771 11943 36777
rect 11885 36768 11897 36771
rect 10928 36740 11897 36768
rect 10928 36728 10934 36740
rect 11885 36737 11897 36740
rect 11931 36768 11943 36771
rect 18138 36768 18144 36780
rect 11931 36740 18144 36768
rect 11931 36737 11943 36740
rect 11885 36731 11943 36737
rect 18138 36728 18144 36740
rect 18196 36728 18202 36780
rect 27154 36768 27160 36780
rect 27067 36740 27160 36768
rect 27154 36728 27160 36740
rect 27212 36768 27218 36780
rect 31128 36777 31156 36808
rect 27801 36771 27859 36777
rect 27801 36768 27813 36771
rect 27212 36740 27813 36768
rect 27212 36728 27218 36740
rect 27801 36737 27813 36740
rect 27847 36737 27859 36771
rect 28905 36771 28963 36777
rect 28905 36768 28917 36771
rect 27801 36731 27859 36737
rect 28368 36740 28917 36768
rect 1854 36632 1860 36644
rect 1815 36604 1860 36632
rect 1854 36592 1860 36604
rect 1912 36592 1918 36644
rect 28368 36576 28396 36740
rect 28905 36737 28917 36740
rect 28951 36737 28963 36771
rect 28905 36731 28963 36737
rect 31113 36771 31171 36777
rect 31113 36737 31125 36771
rect 31159 36737 31171 36771
rect 31312 36768 31340 36867
rect 35526 36864 35532 36876
rect 35584 36864 35590 36916
rect 34885 36839 34943 36845
rect 34885 36805 34897 36839
rect 34931 36836 34943 36839
rect 36265 36839 36323 36845
rect 36265 36836 36277 36839
rect 34931 36808 36277 36836
rect 34931 36805 34943 36808
rect 34885 36799 34943 36805
rect 36265 36805 36277 36808
rect 36311 36836 36323 36839
rect 37366 36836 37372 36848
rect 36311 36808 37372 36836
rect 36311 36805 36323 36808
rect 36265 36799 36323 36805
rect 37366 36796 37372 36808
rect 37424 36796 37430 36848
rect 35345 36771 35403 36777
rect 35345 36768 35357 36771
rect 31312 36740 35357 36768
rect 31113 36731 31171 36737
rect 35345 36737 35357 36740
rect 35391 36737 35403 36771
rect 35345 36731 35403 36737
rect 3234 36564 3240 36576
rect 3195 36536 3240 36564
rect 3234 36524 3240 36536
rect 3292 36524 3298 36576
rect 13909 36567 13967 36573
rect 13909 36533 13921 36567
rect 13955 36564 13967 36567
rect 13998 36564 14004 36576
rect 13955 36536 14004 36564
rect 13955 36533 13967 36536
rect 13909 36527 13967 36533
rect 13998 36524 14004 36536
rect 14056 36524 14062 36576
rect 28350 36564 28356 36576
rect 28311 36536 28356 36564
rect 28350 36524 28356 36536
rect 28408 36524 28414 36576
rect 36170 36564 36176 36576
rect 36131 36536 36176 36564
rect 36170 36524 36176 36536
rect 36228 36524 36234 36576
rect 1104 36474 36892 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 36892 36474
rect 1104 36400 36892 36422
rect 17678 36320 17684 36372
rect 17736 36360 17742 36372
rect 28350 36360 28356 36372
rect 17736 36332 28356 36360
rect 17736 36320 17742 36332
rect 28350 36320 28356 36332
rect 28408 36320 28414 36372
rect 35618 36360 35624 36372
rect 35579 36332 35624 36360
rect 35618 36320 35624 36332
rect 35676 36320 35682 36372
rect 1765 36295 1823 36301
rect 1765 36261 1777 36295
rect 1811 36292 1823 36295
rect 2498 36292 2504 36304
rect 1811 36264 2504 36292
rect 1811 36261 1823 36264
rect 1765 36255 1823 36261
rect 2498 36252 2504 36264
rect 2556 36252 2562 36304
rect 26697 36295 26755 36301
rect 26697 36261 26709 36295
rect 26743 36292 26755 36295
rect 26743 36264 35894 36292
rect 26743 36261 26755 36264
rect 26697 36255 26755 36261
rect 658 36116 664 36168
rect 716 36156 722 36168
rect 1581 36159 1639 36165
rect 1581 36156 1593 36159
rect 716 36128 1593 36156
rect 716 36116 722 36128
rect 1581 36125 1593 36128
rect 1627 36156 1639 36159
rect 2225 36159 2283 36165
rect 2225 36156 2237 36159
rect 1627 36128 2237 36156
rect 1627 36125 1639 36128
rect 1581 36119 1639 36125
rect 2225 36125 2237 36128
rect 2271 36125 2283 36159
rect 2225 36119 2283 36125
rect 26418 36116 26424 36168
rect 26476 36156 26482 36168
rect 26513 36159 26571 36165
rect 26513 36156 26525 36159
rect 26476 36128 26525 36156
rect 26476 36116 26482 36128
rect 26513 36125 26525 36128
rect 26559 36156 26571 36159
rect 27157 36159 27215 36165
rect 27157 36156 27169 36159
rect 26559 36128 27169 36156
rect 26559 36125 26571 36128
rect 26513 36119 26571 36125
rect 27157 36125 27169 36128
rect 27203 36125 27215 36159
rect 35866 36156 35894 36264
rect 36081 36159 36139 36165
rect 36081 36156 36093 36159
rect 35866 36128 36093 36156
rect 27157 36119 27215 36125
rect 36081 36125 36093 36128
rect 36127 36125 36139 36159
rect 36081 36119 36139 36125
rect 36262 36020 36268 36032
rect 36223 35992 36268 36020
rect 36262 35980 36268 35992
rect 36320 35980 36326 36032
rect 1104 35930 36892 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 36892 35930
rect 1104 35856 36892 35878
rect 1578 35612 1584 35624
rect 1539 35584 1584 35612
rect 1578 35572 1584 35584
rect 1636 35572 1642 35624
rect 1857 35615 1915 35621
rect 1857 35581 1869 35615
rect 1903 35612 1915 35615
rect 2682 35612 2688 35624
rect 1903 35584 2688 35612
rect 1903 35581 1915 35584
rect 1857 35575 1915 35581
rect 2682 35572 2688 35584
rect 2740 35572 2746 35624
rect 1104 35386 36892 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 36892 35386
rect 1104 35312 36892 35334
rect 1578 35272 1584 35284
rect 1539 35244 1584 35272
rect 1578 35232 1584 35244
rect 1636 35232 1642 35284
rect 27154 35028 27160 35080
rect 27212 35068 27218 35080
rect 36081 35071 36139 35077
rect 36081 35068 36093 35071
rect 27212 35040 36093 35068
rect 27212 35028 27218 35040
rect 36081 35037 36093 35040
rect 36127 35037 36139 35071
rect 36354 35068 36360 35080
rect 36315 35040 36360 35068
rect 36081 35031 36139 35037
rect 36354 35028 36360 35040
rect 36412 35028 36418 35080
rect 1104 34842 36892 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 36892 34842
rect 1104 34768 36892 34790
rect 36354 34728 36360 34740
rect 36315 34700 36360 34728
rect 36354 34688 36360 34700
rect 36412 34688 36418 34740
rect 1104 34298 36892 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 36892 34298
rect 1104 34224 36892 34246
rect 1104 33754 36892 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 36892 33754
rect 1104 33680 36892 33702
rect 1104 33210 36892 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 36892 33210
rect 1104 33136 36892 33158
rect 18874 33096 18880 33108
rect 18835 33068 18880 33096
rect 18874 33056 18880 33068
rect 18932 33056 18938 33108
rect 18230 32852 18236 32904
rect 18288 32892 18294 32904
rect 18693 32895 18751 32901
rect 18693 32892 18705 32895
rect 18288 32864 18705 32892
rect 18288 32852 18294 32864
rect 18693 32861 18705 32864
rect 18739 32892 18751 32895
rect 19429 32895 19487 32901
rect 19429 32892 19441 32895
rect 18739 32864 19441 32892
rect 18739 32861 18751 32864
rect 18693 32855 18751 32861
rect 19429 32861 19441 32864
rect 19475 32861 19487 32895
rect 19429 32855 19487 32861
rect 24581 32895 24639 32901
rect 24581 32861 24593 32895
rect 24627 32892 24639 32895
rect 25225 32895 25283 32901
rect 25225 32892 25237 32895
rect 24627 32864 25237 32892
rect 24627 32861 24639 32864
rect 24581 32855 24639 32861
rect 25225 32861 25237 32864
rect 25271 32861 25283 32895
rect 25225 32855 25283 32861
rect 13814 32784 13820 32836
rect 13872 32824 13878 32836
rect 24596 32824 24624 32855
rect 13872 32796 24624 32824
rect 24673 32827 24731 32833
rect 13872 32784 13878 32796
rect 24673 32793 24685 32827
rect 24719 32824 24731 32827
rect 31018 32824 31024 32836
rect 24719 32796 31024 32824
rect 24719 32793 24731 32796
rect 24673 32787 24731 32793
rect 31018 32784 31024 32796
rect 31076 32784 31082 32836
rect 35621 32827 35679 32833
rect 35621 32793 35633 32827
rect 35667 32824 35679 32827
rect 36262 32824 36268 32836
rect 35667 32796 36268 32824
rect 35667 32793 35679 32796
rect 35621 32787 35679 32793
rect 36262 32784 36268 32796
rect 36320 32784 36326 32836
rect 36173 32759 36231 32765
rect 36173 32725 36185 32759
rect 36219 32756 36231 32759
rect 36538 32756 36544 32768
rect 36219 32728 36544 32756
rect 36219 32725 36231 32728
rect 36173 32719 36231 32725
rect 36538 32716 36544 32728
rect 36596 32716 36602 32768
rect 1104 32666 36892 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 36892 32666
rect 1104 32592 36892 32614
rect 1578 32348 1584 32360
rect 1539 32320 1584 32348
rect 1578 32308 1584 32320
rect 1636 32308 1642 32360
rect 1857 32351 1915 32357
rect 1857 32317 1869 32351
rect 1903 32348 1915 32351
rect 2774 32348 2780 32360
rect 1903 32320 2780 32348
rect 1903 32317 1915 32320
rect 1857 32311 1915 32317
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 1104 32122 36892 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 36892 32122
rect 1104 32048 36892 32070
rect 1578 32008 1584 32020
rect 1539 31980 1584 32008
rect 1578 31968 1584 31980
rect 1636 31968 1642 32020
rect 10045 32011 10103 32017
rect 10045 31977 10057 32011
rect 10091 32008 10103 32011
rect 10778 32008 10784 32020
rect 10091 31980 10784 32008
rect 10091 31977 10103 31980
rect 10045 31971 10103 31977
rect 10778 31968 10784 31980
rect 10836 31968 10842 32020
rect 35802 31900 35808 31952
rect 35860 31940 35866 31952
rect 36265 31943 36323 31949
rect 36265 31940 36277 31943
rect 35860 31912 36277 31940
rect 35860 31900 35866 31912
rect 36265 31909 36277 31912
rect 36311 31909 36323 31943
rect 36265 31903 36323 31909
rect 5718 31764 5724 31816
rect 5776 31804 5782 31816
rect 9953 31807 10011 31813
rect 9953 31804 9965 31807
rect 5776 31776 9965 31804
rect 5776 31764 5782 31776
rect 9953 31773 9965 31776
rect 9999 31773 10011 31807
rect 10686 31804 10692 31816
rect 10647 31776 10692 31804
rect 9953 31767 10011 31773
rect 10686 31764 10692 31776
rect 10744 31764 10750 31816
rect 10781 31807 10839 31813
rect 10781 31773 10793 31807
rect 10827 31804 10839 31807
rect 10870 31804 10876 31816
rect 10827 31776 10876 31804
rect 10827 31773 10839 31776
rect 10781 31767 10839 31773
rect 10870 31764 10876 31776
rect 10928 31764 10934 31816
rect 27798 31764 27804 31816
rect 27856 31804 27862 31816
rect 36081 31807 36139 31813
rect 36081 31804 36093 31807
rect 27856 31776 36093 31804
rect 27856 31764 27862 31776
rect 36081 31773 36093 31776
rect 36127 31773 36139 31807
rect 36081 31767 36139 31773
rect 1104 31578 36892 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 36892 31578
rect 1104 31504 36892 31526
rect 9398 31424 9404 31476
rect 9456 31464 9462 31476
rect 10321 31467 10379 31473
rect 10321 31464 10333 31467
rect 9456 31436 10333 31464
rect 9456 31424 9462 31436
rect 10321 31433 10333 31436
rect 10367 31433 10379 31467
rect 10321 31427 10379 31433
rect 10413 31331 10471 31337
rect 10413 31297 10425 31331
rect 10459 31328 10471 31331
rect 12894 31328 12900 31340
rect 10459 31300 12900 31328
rect 10459 31297 10471 31300
rect 10413 31291 10471 31297
rect 12894 31288 12900 31300
rect 12952 31288 12958 31340
rect 1104 31034 36892 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 36892 31034
rect 1104 30960 36892 30982
rect 21361 30923 21419 30929
rect 21361 30889 21373 30923
rect 21407 30920 21419 30923
rect 24578 30920 24584 30932
rect 21407 30892 24584 30920
rect 21407 30889 21419 30892
rect 21361 30883 21419 30889
rect 24578 30880 24584 30892
rect 24636 30880 24642 30932
rect 1857 30719 1915 30725
rect 1857 30685 1869 30719
rect 1903 30716 1915 30719
rect 13170 30716 13176 30728
rect 1903 30688 13176 30716
rect 1903 30685 1915 30688
rect 1857 30679 1915 30685
rect 13170 30676 13176 30688
rect 13228 30676 13234 30728
rect 21174 30676 21180 30728
rect 21232 30716 21238 30728
rect 21269 30719 21327 30725
rect 21269 30716 21281 30719
rect 21232 30688 21281 30716
rect 21232 30676 21238 30688
rect 21269 30685 21281 30688
rect 21315 30685 21327 30719
rect 21269 30679 21327 30685
rect 1670 30580 1676 30592
rect 1631 30552 1676 30580
rect 1670 30540 1676 30552
rect 1728 30540 1734 30592
rect 1104 30490 36892 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 36892 30490
rect 1104 30416 36892 30438
rect 13170 30376 13176 30388
rect 13131 30348 13176 30376
rect 13170 30336 13176 30348
rect 13228 30336 13234 30388
rect 2314 30268 2320 30320
rect 2372 30308 2378 30320
rect 4893 30311 4951 30317
rect 4893 30308 4905 30311
rect 2372 30280 4905 30308
rect 2372 30268 2378 30280
rect 4893 30277 4905 30280
rect 4939 30277 4951 30311
rect 4893 30271 4951 30277
rect 4614 30200 4620 30252
rect 4672 30240 4678 30252
rect 4801 30243 4859 30249
rect 4801 30240 4813 30243
rect 4672 30212 4813 30240
rect 4672 30200 4678 30212
rect 4801 30209 4813 30212
rect 4847 30209 4859 30243
rect 4801 30203 4859 30209
rect 12437 30243 12495 30249
rect 12437 30209 12449 30243
rect 12483 30240 12495 30243
rect 12526 30240 12532 30252
rect 12483 30212 12532 30240
rect 12483 30209 12495 30212
rect 12437 30203 12495 30209
rect 12526 30200 12532 30212
rect 12584 30200 12590 30252
rect 12618 30200 12624 30252
rect 12676 30240 12682 30252
rect 13357 30243 13415 30249
rect 13357 30240 13369 30243
rect 12676 30212 13369 30240
rect 12676 30200 12682 30212
rect 13357 30209 13369 30212
rect 13403 30240 13415 30243
rect 22649 30243 22707 30249
rect 13403 30212 13952 30240
rect 13403 30209 13415 30212
rect 13357 30203 13415 30209
rect 12250 30104 12256 30116
rect 12211 30076 12256 30104
rect 12250 30064 12256 30076
rect 12308 30064 12314 30116
rect 13924 30113 13952 30212
rect 22649 30209 22661 30243
rect 22695 30240 22707 30243
rect 27430 30240 27436 30252
rect 22695 30212 27436 30240
rect 22695 30209 22707 30212
rect 22649 30203 22707 30209
rect 27430 30200 27436 30212
rect 27488 30200 27494 30252
rect 13909 30107 13967 30113
rect 13909 30073 13921 30107
rect 13955 30104 13967 30107
rect 32950 30104 32956 30116
rect 13955 30076 32956 30104
rect 13955 30073 13967 30076
rect 13909 30067 13967 30073
rect 32950 30064 32956 30076
rect 33008 30064 33014 30116
rect 22554 30036 22560 30048
rect 22515 30008 22560 30036
rect 22554 29996 22560 30008
rect 22612 29996 22618 30048
rect 1104 29946 36892 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 36892 29946
rect 1104 29872 36892 29894
rect 22189 29631 22247 29637
rect 22189 29597 22201 29631
rect 22235 29628 22247 29631
rect 22741 29631 22799 29637
rect 22741 29628 22753 29631
rect 22235 29600 22753 29628
rect 22235 29597 22247 29600
rect 22189 29591 22247 29597
rect 22741 29597 22753 29600
rect 22787 29628 22799 29631
rect 27154 29628 27160 29640
rect 22787 29600 27160 29628
rect 22787 29597 22799 29600
rect 22741 29591 22799 29597
rect 27154 29588 27160 29600
rect 27212 29588 27218 29640
rect 35621 29563 35679 29569
rect 35621 29529 35633 29563
rect 35667 29560 35679 29563
rect 36262 29560 36268 29572
rect 35667 29532 36268 29560
rect 35667 29529 35679 29532
rect 35621 29523 35679 29529
rect 36262 29520 36268 29532
rect 36320 29520 36326 29572
rect 12526 29492 12532 29504
rect 12487 29464 12532 29492
rect 12526 29452 12532 29464
rect 12584 29452 12590 29504
rect 17218 29452 17224 29504
rect 17276 29492 17282 29504
rect 22097 29495 22155 29501
rect 22097 29492 22109 29495
rect 17276 29464 22109 29492
rect 17276 29452 17282 29464
rect 22097 29461 22109 29464
rect 22143 29461 22155 29495
rect 22097 29455 22155 29461
rect 35986 29452 35992 29504
rect 36044 29492 36050 29504
rect 36173 29495 36231 29501
rect 36173 29492 36185 29495
rect 36044 29464 36185 29492
rect 36044 29452 36050 29464
rect 36173 29461 36185 29464
rect 36219 29461 36231 29495
rect 36173 29455 36231 29461
rect 1104 29402 36892 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 36892 29402
rect 1104 29328 36892 29350
rect 16114 29288 16120 29300
rect 16075 29260 16120 29288
rect 16114 29248 16120 29260
rect 16172 29248 16178 29300
rect 1578 29152 1584 29164
rect 1539 29124 1584 29152
rect 1578 29112 1584 29124
rect 1636 29152 1642 29164
rect 2225 29155 2283 29161
rect 2225 29152 2237 29155
rect 1636 29124 2237 29152
rect 1636 29112 1642 29124
rect 2225 29121 2237 29124
rect 2271 29121 2283 29155
rect 2225 29115 2283 29121
rect 15657 29155 15715 29161
rect 15657 29121 15669 29155
rect 15703 29152 15715 29155
rect 16132 29152 16160 29248
rect 15703 29124 16160 29152
rect 15703 29121 15715 29124
rect 15657 29115 15715 29121
rect 1762 29016 1768 29028
rect 1723 28988 1768 29016
rect 1762 28976 1768 28988
rect 1820 28976 1826 29028
rect 15565 29019 15623 29025
rect 15565 28985 15577 29019
rect 15611 29016 15623 29019
rect 15654 29016 15660 29028
rect 15611 28988 15660 29016
rect 15611 28985 15623 28988
rect 15565 28979 15623 28985
rect 15654 28976 15660 28988
rect 15712 28976 15718 29028
rect 1104 28858 36892 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 36892 28858
rect 1104 28784 36892 28806
rect 14645 28747 14703 28753
rect 14645 28713 14657 28747
rect 14691 28744 14703 28747
rect 16850 28744 16856 28756
rect 14691 28716 16856 28744
rect 14691 28713 14703 28716
rect 14645 28707 14703 28713
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 13906 28500 13912 28552
rect 13964 28540 13970 28552
rect 14461 28543 14519 28549
rect 14461 28540 14473 28543
rect 13964 28512 14473 28540
rect 13964 28500 13970 28512
rect 14461 28509 14473 28512
rect 14507 28540 14519 28543
rect 15105 28543 15163 28549
rect 15105 28540 15117 28543
rect 14507 28512 15117 28540
rect 14507 28509 14519 28512
rect 14461 28503 14519 28509
rect 15105 28509 15117 28512
rect 15151 28509 15163 28543
rect 15105 28503 15163 28509
rect 1104 28314 36892 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 36892 28314
rect 1104 28240 36892 28262
rect 35621 28067 35679 28073
rect 35621 28033 35633 28067
rect 35667 28064 35679 28067
rect 36262 28064 36268 28076
rect 35667 28036 36268 28064
rect 35667 28033 35679 28036
rect 35621 28027 35679 28033
rect 36262 28024 36268 28036
rect 36320 28024 36326 28076
rect 15289 27931 15347 27937
rect 15289 27897 15301 27931
rect 15335 27928 15347 27931
rect 15562 27928 15568 27940
rect 15335 27900 15568 27928
rect 15335 27897 15347 27900
rect 15289 27891 15347 27897
rect 15562 27888 15568 27900
rect 15620 27888 15626 27940
rect 35894 27888 35900 27940
rect 35952 27928 35958 27940
rect 36081 27931 36139 27937
rect 36081 27928 36093 27931
rect 35952 27900 36093 27928
rect 35952 27888 35958 27900
rect 36081 27897 36093 27900
rect 36127 27897 36139 27931
rect 36081 27891 36139 27897
rect 1854 27820 1860 27872
rect 1912 27860 1918 27872
rect 1949 27863 2007 27869
rect 1949 27860 1961 27863
rect 1912 27832 1961 27860
rect 1912 27820 1918 27832
rect 1949 27829 1961 27832
rect 1995 27829 2007 27863
rect 1949 27823 2007 27829
rect 11977 27863 12035 27869
rect 11977 27829 11989 27863
rect 12023 27860 12035 27863
rect 12066 27860 12072 27872
rect 12023 27832 12072 27860
rect 12023 27829 12035 27832
rect 11977 27823 12035 27829
rect 12066 27820 12072 27832
rect 12124 27820 12130 27872
rect 15470 27820 15476 27872
rect 15528 27860 15534 27872
rect 15749 27863 15807 27869
rect 15749 27860 15761 27863
rect 15528 27832 15761 27860
rect 15528 27820 15534 27832
rect 15749 27829 15761 27832
rect 15795 27829 15807 27863
rect 15749 27823 15807 27829
rect 1104 27770 36892 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 36892 27770
rect 1104 27696 36892 27718
rect 12618 27588 12624 27600
rect 12579 27560 12624 27588
rect 12618 27548 12624 27560
rect 12676 27548 12682 27600
rect 1854 27452 1860 27464
rect 1815 27424 1860 27452
rect 1854 27412 1860 27424
rect 1912 27412 1918 27464
rect 2498 27452 2504 27464
rect 2459 27424 2504 27452
rect 2498 27412 2504 27424
rect 2556 27412 2562 27464
rect 15470 27412 15476 27464
rect 15528 27452 15534 27464
rect 15565 27455 15623 27461
rect 15565 27452 15577 27455
rect 15528 27424 15577 27452
rect 15528 27412 15534 27424
rect 15565 27421 15577 27424
rect 15611 27421 15623 27455
rect 15565 27415 15623 27421
rect 2682 27344 2688 27396
rect 2740 27384 2746 27396
rect 16025 27387 16083 27393
rect 16025 27384 16037 27387
rect 2740 27356 16037 27384
rect 2740 27344 2746 27356
rect 16025 27353 16037 27356
rect 16071 27384 16083 27387
rect 16390 27384 16396 27396
rect 16071 27356 16396 27384
rect 16071 27353 16083 27356
rect 16025 27347 16083 27353
rect 16390 27344 16396 27356
rect 16448 27344 16454 27396
rect 1670 27316 1676 27328
rect 1631 27288 1676 27316
rect 1670 27276 1676 27288
rect 1728 27276 1734 27328
rect 2314 27316 2320 27328
rect 2275 27288 2320 27316
rect 2314 27276 2320 27288
rect 2372 27276 2378 27328
rect 10873 27319 10931 27325
rect 10873 27285 10885 27319
rect 10919 27316 10931 27319
rect 11146 27316 11152 27328
rect 10919 27288 11152 27316
rect 10919 27285 10931 27288
rect 10873 27279 10931 27285
rect 11146 27276 11152 27288
rect 11204 27276 11210 27328
rect 11701 27319 11759 27325
rect 11701 27285 11713 27319
rect 11747 27316 11759 27319
rect 11790 27316 11796 27328
rect 11747 27288 11796 27316
rect 11747 27285 11759 27288
rect 11701 27279 11759 27285
rect 11790 27276 11796 27288
rect 11848 27276 11854 27328
rect 14369 27319 14427 27325
rect 14369 27285 14381 27319
rect 14415 27316 14427 27319
rect 14458 27316 14464 27328
rect 14415 27288 14464 27316
rect 14415 27285 14427 27288
rect 14369 27279 14427 27285
rect 14458 27276 14464 27288
rect 14516 27276 14522 27328
rect 14826 27316 14832 27328
rect 14787 27288 14832 27316
rect 14826 27276 14832 27288
rect 14884 27276 14890 27328
rect 14918 27276 14924 27328
rect 14976 27316 14982 27328
rect 15473 27319 15531 27325
rect 15473 27316 15485 27319
rect 14976 27288 15485 27316
rect 14976 27276 14982 27288
rect 15473 27285 15485 27288
rect 15519 27285 15531 27319
rect 15473 27279 15531 27285
rect 1104 27226 36892 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 36892 27226
rect 1104 27152 36892 27174
rect 5902 27072 5908 27124
rect 5960 27112 5966 27124
rect 5960 27084 13124 27112
rect 5960 27072 5966 27084
rect 8021 27047 8079 27053
rect 8021 27013 8033 27047
rect 8067 27044 8079 27047
rect 8570 27044 8576 27056
rect 8067 27016 8576 27044
rect 8067 27013 8079 27016
rect 8021 27007 8079 27013
rect 8570 27004 8576 27016
rect 8628 27004 8634 27056
rect 11790 27044 11796 27056
rect 11751 27016 11796 27044
rect 11790 27004 11796 27016
rect 11848 27004 11854 27056
rect 11882 27004 11888 27056
rect 11940 27044 11946 27056
rect 13096 27053 13124 27084
rect 13081 27047 13139 27053
rect 11940 27016 11985 27044
rect 11940 27004 11946 27016
rect 13081 27013 13093 27047
rect 13127 27013 13139 27047
rect 13081 27007 13139 27013
rect 13633 27047 13691 27053
rect 13633 27013 13645 27047
rect 13679 27044 13691 27047
rect 13814 27044 13820 27056
rect 13679 27016 13820 27044
rect 13679 27013 13691 27016
rect 13633 27007 13691 27013
rect 13814 27004 13820 27016
rect 13872 27044 13878 27056
rect 14182 27044 14188 27056
rect 13872 27016 14188 27044
rect 13872 27004 13878 27016
rect 14182 27004 14188 27016
rect 14240 27004 14246 27056
rect 14918 27044 14924 27056
rect 14879 27016 14924 27044
rect 14918 27004 14924 27016
rect 14976 27004 14982 27056
rect 15013 27047 15071 27053
rect 15013 27013 15025 27047
rect 15059 27044 15071 27047
rect 15654 27044 15660 27056
rect 15059 27016 15660 27044
rect 15059 27013 15071 27016
rect 15013 27007 15071 27013
rect 15654 27004 15660 27016
rect 15712 27004 15718 27056
rect 15749 27047 15807 27053
rect 15749 27013 15761 27047
rect 15795 27044 15807 27047
rect 16666 27044 16672 27056
rect 15795 27016 16672 27044
rect 15795 27013 15807 27016
rect 15749 27007 15807 27013
rect 16666 27004 16672 27016
rect 16724 27004 16730 27056
rect 2133 26979 2191 26985
rect 2133 26945 2145 26979
rect 2179 26976 2191 26979
rect 2777 26979 2835 26985
rect 2777 26976 2789 26979
rect 2179 26948 2789 26976
rect 2179 26945 2191 26948
rect 2133 26939 2191 26945
rect 2777 26945 2789 26948
rect 2823 26976 2835 26979
rect 2958 26976 2964 26988
rect 2823 26948 2964 26976
rect 2823 26945 2835 26948
rect 2777 26939 2835 26945
rect 2958 26936 2964 26948
rect 3016 26936 3022 26988
rect 11146 26976 11152 26988
rect 11059 26948 11152 26976
rect 11146 26936 11152 26948
rect 11204 26936 11210 26988
rect 16390 26936 16396 26988
rect 16448 26976 16454 26988
rect 17037 26979 17095 26985
rect 17037 26976 17049 26979
rect 16448 26948 17049 26976
rect 16448 26936 16454 26948
rect 17037 26945 17049 26948
rect 17083 26976 17095 26979
rect 17497 26979 17555 26985
rect 17497 26976 17509 26979
rect 17083 26948 17509 26976
rect 17083 26945 17095 26948
rect 17037 26939 17095 26945
rect 17497 26945 17509 26948
rect 17543 26945 17555 26979
rect 17497 26939 17555 26945
rect 7926 26908 7932 26920
rect 7887 26880 7932 26908
rect 7926 26868 7932 26880
rect 7984 26868 7990 26920
rect 11164 26908 11192 26936
rect 12066 26908 12072 26920
rect 11164 26880 12072 26908
rect 12066 26868 12072 26880
rect 12124 26868 12130 26920
rect 12437 26911 12495 26917
rect 12437 26877 12449 26911
rect 12483 26908 12495 26911
rect 12989 26911 13047 26917
rect 12989 26908 13001 26911
rect 12483 26880 13001 26908
rect 12483 26877 12495 26880
rect 12437 26871 12495 26877
rect 12989 26877 13001 26880
rect 13035 26877 13047 26911
rect 12989 26871 13047 26877
rect 14737 26911 14795 26917
rect 14737 26877 14749 26911
rect 14783 26908 14795 26911
rect 15838 26908 15844 26920
rect 14783 26880 15844 26908
rect 14783 26877 14795 26880
rect 14737 26871 14795 26877
rect 1486 26800 1492 26852
rect 1544 26840 1550 26852
rect 2593 26843 2651 26849
rect 2593 26840 2605 26843
rect 1544 26812 2605 26840
rect 1544 26800 1550 26812
rect 2593 26809 2605 26812
rect 2639 26809 2651 26843
rect 2593 26803 2651 26809
rect 4982 26800 4988 26852
rect 5040 26840 5046 26852
rect 8481 26843 8539 26849
rect 8481 26840 8493 26843
rect 5040 26812 8493 26840
rect 5040 26800 5046 26812
rect 8481 26809 8493 26812
rect 8527 26840 8539 26843
rect 9214 26840 9220 26852
rect 8527 26812 9220 26840
rect 8527 26809 8539 26812
rect 8481 26803 8539 26809
rect 9214 26800 9220 26812
rect 9272 26800 9278 26852
rect 10594 26800 10600 26852
rect 10652 26840 10658 26852
rect 12452 26840 12480 26871
rect 15838 26868 15844 26880
rect 15896 26868 15902 26920
rect 16301 26911 16359 26917
rect 16301 26877 16313 26911
rect 16347 26908 16359 26911
rect 17586 26908 17592 26920
rect 16347 26880 17592 26908
rect 16347 26877 16359 26880
rect 16301 26871 16359 26877
rect 17586 26868 17592 26880
rect 17644 26868 17650 26920
rect 10652 26812 12480 26840
rect 10652 26800 10658 26812
rect 1946 26732 1952 26784
rect 2004 26772 2010 26784
rect 2041 26775 2099 26781
rect 2041 26772 2053 26775
rect 2004 26744 2053 26772
rect 2004 26732 2010 26744
rect 2041 26741 2053 26744
rect 2087 26741 2099 26775
rect 10502 26772 10508 26784
rect 10463 26744 10508 26772
rect 2041 26735 2099 26741
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 10962 26732 10968 26784
rect 11020 26772 11026 26784
rect 11057 26775 11115 26781
rect 11057 26772 11069 26775
rect 11020 26744 11069 26772
rect 11020 26732 11026 26744
rect 11057 26741 11069 26744
rect 11103 26741 11115 26775
rect 11057 26735 11115 26741
rect 16574 26732 16580 26784
rect 16632 26772 16638 26784
rect 16945 26775 17003 26781
rect 16945 26772 16957 26775
rect 16632 26744 16957 26772
rect 16632 26732 16638 26744
rect 16945 26741 16957 26744
rect 16991 26741 17003 26775
rect 16945 26735 17003 26741
rect 1104 26682 36892 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 36892 26682
rect 1104 26608 36892 26630
rect 6730 26528 6736 26580
rect 6788 26568 6794 26580
rect 11701 26571 11759 26577
rect 6788 26540 11192 26568
rect 6788 26528 6794 26540
rect 1673 26503 1731 26509
rect 1673 26469 1685 26503
rect 1719 26500 1731 26503
rect 1854 26500 1860 26512
rect 1719 26472 1860 26500
rect 1719 26469 1731 26472
rect 1673 26463 1731 26469
rect 1854 26460 1860 26472
rect 1912 26460 1918 26512
rect 8202 26460 8208 26512
rect 8260 26500 8266 26512
rect 10505 26503 10563 26509
rect 10505 26500 10517 26503
rect 8260 26472 10517 26500
rect 8260 26460 8266 26472
rect 10505 26469 10517 26472
rect 10551 26500 10563 26503
rect 10594 26500 10600 26512
rect 10551 26472 10600 26500
rect 10551 26469 10563 26472
rect 10505 26463 10563 26469
rect 10594 26460 10600 26472
rect 10652 26460 10658 26512
rect 2409 26435 2467 26441
rect 2409 26401 2421 26435
rect 2455 26432 2467 26435
rect 5258 26432 5264 26444
rect 2455 26404 5264 26432
rect 2455 26401 2467 26404
rect 2409 26395 2467 26401
rect 5258 26392 5264 26404
rect 5316 26392 5322 26444
rect 7926 26432 7932 26444
rect 7887 26404 7932 26432
rect 7926 26392 7932 26404
rect 7984 26392 7990 26444
rect 9214 26432 9220 26444
rect 9175 26404 9220 26432
rect 9214 26392 9220 26404
rect 9272 26392 9278 26444
rect 9861 26435 9919 26441
rect 9861 26401 9873 26435
rect 9907 26432 9919 26435
rect 10686 26432 10692 26444
rect 9907 26404 10692 26432
rect 9907 26401 9919 26404
rect 9861 26395 9919 26401
rect 10686 26392 10692 26404
rect 10744 26432 10750 26444
rect 11057 26435 11115 26441
rect 11057 26432 11069 26435
rect 10744 26404 11069 26432
rect 10744 26392 10750 26404
rect 11057 26401 11069 26404
rect 11103 26401 11115 26435
rect 11164 26432 11192 26540
rect 11701 26537 11713 26571
rect 11747 26568 11759 26571
rect 11882 26568 11888 26580
rect 11747 26540 11888 26568
rect 11747 26537 11759 26540
rect 11701 26531 11759 26537
rect 11882 26528 11888 26540
rect 11940 26528 11946 26580
rect 17218 26568 17224 26580
rect 16546 26540 17224 26568
rect 12345 26503 12403 26509
rect 12345 26469 12357 26503
rect 12391 26500 12403 26503
rect 12434 26500 12440 26512
rect 12391 26472 12440 26500
rect 12391 26469 12403 26472
rect 12345 26463 12403 26469
rect 12434 26460 12440 26472
rect 12492 26460 12498 26512
rect 11164 26404 12848 26432
rect 11057 26395 11115 26401
rect 1670 26324 1676 26376
rect 1728 26364 1734 26376
rect 1857 26367 1915 26373
rect 1857 26364 1869 26367
rect 1728 26336 1869 26364
rect 1728 26324 1734 26336
rect 1857 26333 1869 26336
rect 1903 26333 1915 26367
rect 1857 26327 1915 26333
rect 2501 26367 2559 26373
rect 2501 26333 2513 26367
rect 2547 26364 2559 26367
rect 3602 26364 3608 26376
rect 2547 26336 3608 26364
rect 2547 26333 2559 26336
rect 2501 26327 2559 26333
rect 3602 26324 3608 26336
rect 3660 26324 3666 26376
rect 11609 26367 11667 26373
rect 11609 26333 11621 26367
rect 11655 26364 11667 26367
rect 12250 26364 12256 26376
rect 11655 26336 12256 26364
rect 11655 26333 11667 26336
rect 11609 26327 11667 26333
rect 12250 26324 12256 26336
rect 12308 26324 12314 26376
rect 12437 26367 12495 26373
rect 12437 26333 12449 26367
rect 12483 26364 12495 26367
rect 12618 26364 12624 26376
rect 12483 26336 12624 26364
rect 12483 26333 12495 26336
rect 12437 26327 12495 26333
rect 12618 26324 12624 26336
rect 12676 26324 12682 26376
rect 2682 26256 2688 26308
rect 2740 26296 2746 26308
rect 2961 26299 3019 26305
rect 2961 26296 2973 26299
rect 2740 26268 2973 26296
rect 2740 26256 2746 26268
rect 2961 26265 2973 26268
rect 3007 26265 3019 26299
rect 9766 26296 9772 26308
rect 9727 26268 9772 26296
rect 2961 26259 3019 26265
rect 9766 26256 9772 26268
rect 9824 26256 9830 26308
rect 10962 26296 10968 26308
rect 10923 26268 10968 26296
rect 10962 26256 10968 26268
rect 11020 26256 11026 26308
rect 12820 26228 12848 26404
rect 12894 26392 12900 26444
rect 12952 26432 12958 26444
rect 13541 26435 13599 26441
rect 12952 26404 12997 26432
rect 12952 26392 12958 26404
rect 13541 26401 13553 26435
rect 13587 26432 13599 26435
rect 15838 26432 15844 26444
rect 13587 26404 15844 26432
rect 13587 26401 13599 26404
rect 13541 26395 13599 26401
rect 15838 26392 15844 26404
rect 15896 26392 15902 26444
rect 16025 26435 16083 26441
rect 16025 26401 16037 26435
rect 16071 26432 16083 26435
rect 16546 26432 16574 26540
rect 17218 26528 17224 26540
rect 17276 26528 17282 26580
rect 17494 26500 17500 26512
rect 16684 26472 17500 26500
rect 16684 26441 16712 26472
rect 17494 26460 17500 26472
rect 17552 26460 17558 26512
rect 35802 26460 35808 26512
rect 35860 26500 35866 26512
rect 36265 26503 36323 26509
rect 36265 26500 36277 26503
rect 35860 26472 36277 26500
rect 35860 26460 35866 26472
rect 36265 26469 36277 26472
rect 36311 26469 36323 26503
rect 36265 26463 36323 26469
rect 16071 26404 16574 26432
rect 16669 26435 16727 26441
rect 16071 26401 16083 26404
rect 16025 26395 16083 26401
rect 16669 26401 16681 26435
rect 16715 26401 16727 26435
rect 17310 26432 17316 26444
rect 17271 26404 17316 26432
rect 16669 26395 16727 26401
rect 17310 26392 17316 26404
rect 17368 26392 17374 26444
rect 18785 26435 18843 26441
rect 18785 26401 18797 26435
rect 18831 26432 18843 26435
rect 22554 26432 22560 26444
rect 18831 26404 22560 26432
rect 18831 26401 18843 26404
rect 18785 26395 18843 26401
rect 22554 26392 22560 26404
rect 22612 26392 22618 26444
rect 14550 26324 14556 26376
rect 14608 26364 14614 26376
rect 14921 26367 14979 26373
rect 14921 26364 14933 26367
rect 14608 26336 14933 26364
rect 14608 26324 14614 26336
rect 14921 26333 14933 26336
rect 14967 26364 14979 26367
rect 15286 26364 15292 26376
rect 14967 26336 15292 26364
rect 14967 26333 14979 26336
rect 14921 26327 14979 26333
rect 15286 26324 15292 26336
rect 15344 26324 15350 26376
rect 36078 26364 36084 26376
rect 36039 26336 36084 26364
rect 36078 26324 36084 26336
rect 36136 26324 36142 26376
rect 13449 26299 13507 26305
rect 13449 26296 13461 26299
rect 13004 26268 13461 26296
rect 13004 26228 13032 26268
rect 13449 26265 13461 26268
rect 13495 26265 13507 26299
rect 15378 26296 15384 26308
rect 15339 26268 15384 26296
rect 13449 26259 13507 26265
rect 15378 26256 15384 26268
rect 15436 26256 15442 26308
rect 15933 26299 15991 26305
rect 15933 26265 15945 26299
rect 15979 26296 15991 26299
rect 16761 26299 16819 26305
rect 15979 26268 16620 26296
rect 15979 26265 15991 26268
rect 15933 26259 15991 26265
rect 12820 26200 13032 26228
rect 14366 26188 14372 26240
rect 14424 26228 14430 26240
rect 14829 26231 14887 26237
rect 14829 26228 14841 26231
rect 14424 26200 14841 26228
rect 14424 26188 14430 26200
rect 14829 26197 14841 26200
rect 14875 26197 14887 26231
rect 16592 26228 16620 26268
rect 16761 26265 16773 26299
rect 16807 26296 16819 26299
rect 16807 26268 16988 26296
rect 16807 26265 16819 26268
rect 16761 26259 16819 26265
rect 16960 26240 16988 26268
rect 17586 26256 17592 26308
rect 17644 26296 17650 26308
rect 18141 26299 18199 26305
rect 18141 26296 18153 26299
rect 17644 26268 18153 26296
rect 17644 26256 17650 26268
rect 18141 26265 18153 26268
rect 18187 26265 18199 26299
rect 18141 26259 18199 26265
rect 18506 26256 18512 26308
rect 18564 26296 18570 26308
rect 18693 26299 18751 26305
rect 18693 26296 18705 26299
rect 18564 26268 18705 26296
rect 18564 26256 18570 26268
rect 18693 26265 18705 26268
rect 18739 26265 18751 26299
rect 18693 26259 18751 26265
rect 16850 26228 16856 26240
rect 16592 26200 16856 26228
rect 14829 26191 14887 26197
rect 16850 26188 16856 26200
rect 16908 26188 16914 26240
rect 16942 26188 16948 26240
rect 17000 26188 17006 26240
rect 1104 26138 36892 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 36892 26138
rect 1104 26064 36892 26086
rect 3234 25984 3240 26036
rect 3292 26024 3298 26036
rect 8294 26024 8300 26036
rect 3292 25996 8300 26024
rect 3292 25984 3298 25996
rect 8294 25984 8300 25996
rect 8352 25984 8358 26036
rect 8570 26024 8576 26036
rect 8531 25996 8576 26024
rect 8570 25984 8576 25996
rect 8628 25984 8634 26036
rect 9309 26027 9367 26033
rect 9309 25993 9321 26027
rect 9355 26024 9367 26027
rect 9766 26024 9772 26036
rect 9355 25996 9772 26024
rect 9355 25993 9367 25996
rect 9309 25987 9367 25993
rect 9766 25984 9772 25996
rect 9824 25984 9830 26036
rect 15010 26024 15016 26036
rect 12406 25996 15016 26024
rect 2130 25956 2136 25968
rect 2091 25928 2136 25956
rect 2130 25916 2136 25928
rect 2188 25916 2194 25968
rect 2498 25916 2504 25968
rect 2556 25956 2562 25968
rect 5258 25956 5264 25968
rect 2556 25928 3464 25956
rect 5219 25928 5264 25956
rect 2556 25916 2562 25928
rect 2590 25848 2596 25900
rect 2648 25888 2654 25900
rect 3436 25897 3464 25928
rect 5258 25916 5264 25928
rect 5316 25916 5322 25968
rect 9674 25916 9680 25968
rect 9732 25956 9738 25968
rect 10686 25956 10692 25968
rect 9732 25928 10692 25956
rect 9732 25916 9738 25928
rect 10686 25916 10692 25928
rect 10744 25956 10750 25968
rect 12406 25956 12434 25996
rect 15010 25984 15016 25996
rect 15068 25984 15074 26036
rect 17494 26024 17500 26036
rect 16546 25996 17500 26024
rect 13262 25956 13268 25968
rect 10744 25928 12434 25956
rect 13223 25928 13268 25956
rect 10744 25916 10750 25928
rect 13262 25916 13268 25928
rect 13320 25916 13326 25968
rect 14366 25956 14372 25968
rect 14327 25928 14372 25956
rect 14366 25916 14372 25928
rect 14424 25916 14430 25968
rect 14921 25959 14979 25965
rect 14921 25925 14933 25959
rect 14967 25956 14979 25959
rect 16546 25956 16574 25996
rect 17494 25984 17500 25996
rect 17552 25984 17558 26036
rect 14967 25928 16574 25956
rect 14967 25925 14979 25928
rect 14921 25919 14979 25925
rect 17034 25916 17040 25968
rect 17092 25956 17098 25968
rect 17405 25959 17463 25965
rect 17405 25956 17417 25959
rect 17092 25928 17417 25956
rect 17092 25916 17098 25928
rect 17405 25925 17417 25928
rect 17451 25925 17463 25959
rect 17405 25919 17463 25925
rect 2777 25891 2835 25897
rect 2777 25888 2789 25891
rect 2648 25860 2789 25888
rect 2648 25848 2654 25860
rect 2777 25857 2789 25860
rect 2823 25857 2835 25891
rect 2777 25851 2835 25857
rect 3421 25891 3479 25897
rect 3421 25857 3433 25891
rect 3467 25857 3479 25891
rect 3421 25851 3479 25857
rect 8665 25891 8723 25897
rect 8665 25857 8677 25891
rect 8711 25888 8723 25891
rect 8754 25888 8760 25900
rect 8711 25860 8760 25888
rect 8711 25857 8723 25860
rect 8665 25851 8723 25857
rect 8754 25848 8760 25860
rect 8812 25848 8818 25900
rect 9214 25888 9220 25900
rect 9175 25860 9220 25888
rect 9214 25848 9220 25860
rect 9272 25888 9278 25900
rect 9861 25891 9919 25897
rect 9861 25888 9873 25891
rect 9272 25860 9873 25888
rect 9272 25848 9278 25860
rect 9861 25857 9873 25860
rect 9907 25857 9919 25891
rect 9861 25851 9919 25857
rect 10965 25891 11023 25897
rect 10965 25857 10977 25891
rect 11011 25857 11023 25891
rect 12066 25888 12072 25900
rect 12027 25860 12072 25888
rect 10965 25851 11023 25857
rect 1949 25823 2007 25829
rect 1949 25789 1961 25823
rect 1995 25820 2007 25823
rect 2038 25820 2044 25832
rect 1995 25792 2044 25820
rect 1995 25789 2007 25792
rect 1949 25783 2007 25789
rect 2038 25780 2044 25792
rect 2096 25780 2102 25832
rect 2225 25823 2283 25829
rect 2225 25789 2237 25823
rect 2271 25820 2283 25823
rect 2498 25820 2504 25832
rect 2271 25792 2504 25820
rect 2271 25789 2283 25792
rect 2225 25783 2283 25789
rect 2498 25780 2504 25792
rect 2556 25820 2562 25832
rect 2682 25820 2688 25832
rect 2556 25792 2688 25820
rect 2556 25780 2562 25792
rect 2682 25780 2688 25792
rect 2740 25780 2746 25832
rect 4982 25780 4988 25832
rect 5040 25820 5046 25832
rect 5169 25823 5227 25829
rect 5169 25820 5181 25823
rect 5040 25792 5181 25820
rect 5040 25780 5046 25792
rect 5169 25789 5181 25792
rect 5215 25789 5227 25823
rect 5169 25783 5227 25789
rect 7193 25823 7251 25829
rect 7193 25789 7205 25823
rect 7239 25820 7251 25823
rect 10134 25820 10140 25832
rect 7239 25792 10140 25820
rect 7239 25789 7251 25792
rect 7193 25783 7251 25789
rect 10134 25780 10140 25792
rect 10192 25820 10198 25832
rect 10502 25820 10508 25832
rect 10192 25792 10508 25820
rect 10192 25780 10198 25792
rect 10502 25780 10508 25792
rect 10560 25820 10566 25832
rect 10980 25820 11008 25851
rect 12066 25848 12072 25860
rect 12124 25848 12130 25900
rect 15562 25888 15568 25900
rect 15523 25860 15568 25888
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 16025 25891 16083 25897
rect 16025 25857 16037 25891
rect 16071 25857 16083 25891
rect 18230 25888 18236 25900
rect 18143 25860 18236 25888
rect 16025 25851 16083 25857
rect 12710 25820 12716 25832
rect 10560 25792 11008 25820
rect 12671 25792 12716 25820
rect 10560 25780 10566 25792
rect 12710 25780 12716 25792
rect 12768 25780 12774 25832
rect 13354 25820 13360 25832
rect 13315 25792 13360 25820
rect 13354 25780 13360 25792
rect 13412 25780 13418 25832
rect 14277 25823 14335 25829
rect 14277 25789 14289 25823
rect 14323 25789 14335 25823
rect 14277 25783 14335 25789
rect 2869 25755 2927 25761
rect 2869 25721 2881 25755
rect 2915 25752 2927 25755
rect 5718 25752 5724 25764
rect 2915 25724 5580 25752
rect 5679 25724 5724 25752
rect 2915 25721 2927 25724
rect 2869 25715 2927 25721
rect 3510 25684 3516 25696
rect 3471 25656 3516 25684
rect 3510 25644 3516 25656
rect 3568 25644 3574 25696
rect 5552 25684 5580 25724
rect 5718 25712 5724 25724
rect 5776 25712 5782 25764
rect 11330 25712 11336 25764
rect 11388 25752 11394 25764
rect 14292 25752 14320 25783
rect 15286 25780 15292 25832
rect 15344 25820 15350 25832
rect 16040 25820 16068 25851
rect 18230 25848 18236 25860
rect 18288 25888 18294 25900
rect 18785 25891 18843 25897
rect 18785 25888 18797 25891
rect 18288 25860 18797 25888
rect 18288 25848 18294 25860
rect 18785 25857 18797 25860
rect 18831 25888 18843 25891
rect 35894 25888 35900 25900
rect 18831 25860 35900 25888
rect 18831 25857 18843 25860
rect 18785 25851 18843 25857
rect 35894 25848 35900 25860
rect 35952 25848 35958 25900
rect 16574 25820 16580 25832
rect 15344 25792 16068 25820
rect 16132 25792 16580 25820
rect 15344 25780 15350 25792
rect 16132 25752 16160 25792
rect 16574 25780 16580 25792
rect 16632 25780 16638 25832
rect 17218 25780 17224 25832
rect 17276 25820 17282 25832
rect 17494 25820 17500 25832
rect 17276 25792 17500 25820
rect 17276 25780 17282 25792
rect 17494 25780 17500 25792
rect 17552 25780 17558 25832
rect 11388 25724 16160 25752
rect 11388 25712 11394 25724
rect 16206 25712 16212 25764
rect 16264 25752 16270 25764
rect 16945 25755 17003 25761
rect 16945 25752 16957 25755
rect 16264 25724 16957 25752
rect 16264 25712 16270 25724
rect 16945 25721 16957 25724
rect 16991 25721 17003 25755
rect 16945 25715 17003 25721
rect 6822 25684 6828 25696
rect 5552 25656 6828 25684
rect 6822 25644 6828 25656
rect 6880 25644 6886 25696
rect 7926 25684 7932 25696
rect 7887 25656 7932 25684
rect 7926 25644 7932 25656
rect 7984 25644 7990 25696
rect 9953 25687 10011 25693
rect 9953 25653 9965 25687
rect 9999 25684 10011 25687
rect 10502 25684 10508 25696
rect 9999 25656 10508 25684
rect 9999 25653 10011 25656
rect 9953 25647 10011 25653
rect 10502 25644 10508 25656
rect 10560 25644 10566 25696
rect 11057 25687 11115 25693
rect 11057 25653 11069 25687
rect 11103 25684 11115 25687
rect 11238 25684 11244 25696
rect 11103 25656 11244 25684
rect 11103 25653 11115 25656
rect 11057 25647 11115 25653
rect 11238 25644 11244 25656
rect 11296 25644 11302 25696
rect 12158 25684 12164 25696
rect 12119 25656 12164 25684
rect 12158 25644 12164 25656
rect 12216 25644 12222 25696
rect 13814 25644 13820 25696
rect 13872 25684 13878 25696
rect 15473 25687 15531 25693
rect 15473 25684 15485 25687
rect 13872 25656 15485 25684
rect 13872 25644 13878 25656
rect 15473 25653 15485 25656
rect 15519 25653 15531 25687
rect 15473 25647 15531 25653
rect 16117 25687 16175 25693
rect 16117 25653 16129 25687
rect 16163 25684 16175 25687
rect 17770 25684 17776 25696
rect 16163 25656 17776 25684
rect 16163 25653 16175 25656
rect 16117 25647 16175 25653
rect 17770 25644 17776 25656
rect 17828 25644 17834 25696
rect 18138 25684 18144 25696
rect 18099 25656 18144 25684
rect 18138 25644 18144 25656
rect 18196 25644 18202 25696
rect 1104 25594 36892 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 36892 25594
rect 1104 25520 36892 25542
rect 3510 25440 3516 25492
rect 3568 25480 3574 25492
rect 12526 25480 12532 25492
rect 3568 25452 12532 25480
rect 3568 25440 3574 25452
rect 12526 25440 12532 25452
rect 12584 25440 12590 25492
rect 14734 25440 14740 25492
rect 14792 25480 14798 25492
rect 16206 25480 16212 25492
rect 14792 25452 16212 25480
rect 14792 25440 14798 25452
rect 16206 25440 16212 25452
rect 16264 25440 16270 25492
rect 17034 25480 17040 25492
rect 16995 25452 17040 25480
rect 17034 25440 17040 25452
rect 17092 25440 17098 25492
rect 20070 25480 20076 25492
rect 17788 25452 20076 25480
rect 4614 25412 4620 25424
rect 2746 25384 4620 25412
rect 2038 25304 2044 25356
rect 2096 25344 2102 25356
rect 2225 25347 2283 25353
rect 2225 25344 2237 25347
rect 2096 25316 2237 25344
rect 2096 25304 2102 25316
rect 2225 25313 2237 25316
rect 2271 25344 2283 25347
rect 2746 25344 2774 25384
rect 4614 25372 4620 25384
rect 4672 25372 4678 25424
rect 6273 25415 6331 25421
rect 6273 25381 6285 25415
rect 6319 25412 6331 25415
rect 8202 25412 8208 25424
rect 6319 25384 8208 25412
rect 6319 25381 6331 25384
rect 6273 25375 6331 25381
rect 8202 25372 8208 25384
rect 8260 25372 8266 25424
rect 8294 25372 8300 25424
rect 8352 25412 8358 25424
rect 8352 25384 12434 25412
rect 8352 25372 8358 25384
rect 4065 25347 4123 25353
rect 4065 25344 4077 25347
rect 2271 25316 2774 25344
rect 3160 25316 4077 25344
rect 2271 25313 2283 25316
rect 2225 25307 2283 25313
rect 2406 25208 2412 25220
rect 2367 25180 2412 25208
rect 2406 25168 2412 25180
rect 2464 25168 2470 25220
rect 2501 25211 2559 25217
rect 2501 25177 2513 25211
rect 2547 25208 2559 25211
rect 3160 25208 3188 25316
rect 4065 25313 4077 25316
rect 4111 25344 4123 25347
rect 10962 25344 10968 25356
rect 4111 25316 10968 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 10962 25304 10968 25316
rect 11020 25304 11026 25356
rect 11330 25344 11336 25356
rect 11291 25316 11336 25344
rect 11330 25304 11336 25316
rect 11388 25304 11394 25356
rect 12158 25304 12164 25356
rect 12216 25344 12222 25356
rect 12253 25347 12311 25353
rect 12253 25344 12265 25347
rect 12216 25316 12265 25344
rect 12216 25304 12222 25316
rect 12253 25313 12265 25316
rect 12299 25313 12311 25347
rect 12406 25344 12434 25384
rect 13354 25372 13360 25424
rect 13412 25412 13418 25424
rect 17788 25412 17816 25452
rect 20070 25440 20076 25452
rect 20128 25480 20134 25492
rect 20128 25452 20392 25480
rect 20128 25440 20134 25452
rect 13412 25384 17816 25412
rect 13412 25372 13418 25384
rect 17862 25372 17868 25424
rect 17920 25412 17926 25424
rect 20364 25421 20392 25452
rect 18233 25415 18291 25421
rect 18233 25412 18245 25415
rect 17920 25384 18245 25412
rect 17920 25372 17926 25384
rect 18233 25381 18245 25384
rect 18279 25381 18291 25415
rect 18233 25375 18291 25381
rect 20349 25415 20407 25421
rect 20349 25381 20361 25415
rect 20395 25381 20407 25415
rect 20349 25375 20407 25381
rect 14277 25347 14335 25353
rect 14277 25344 14289 25347
rect 12406 25316 14289 25344
rect 12253 25307 12311 25313
rect 14277 25313 14289 25316
rect 14323 25313 14335 25347
rect 14277 25307 14335 25313
rect 17681 25347 17739 25353
rect 17681 25313 17693 25347
rect 17727 25344 17739 25347
rect 18138 25344 18144 25356
rect 17727 25316 18144 25344
rect 17727 25313 17739 25316
rect 17681 25307 17739 25313
rect 18138 25304 18144 25316
rect 18196 25304 18202 25356
rect 20901 25347 20959 25353
rect 20901 25313 20913 25347
rect 20947 25344 20959 25347
rect 22554 25344 22560 25356
rect 20947 25316 22560 25344
rect 20947 25313 20959 25316
rect 20901 25307 20959 25313
rect 22554 25304 22560 25316
rect 22612 25304 22618 25356
rect 3326 25276 3332 25288
rect 3287 25248 3332 25276
rect 3326 25236 3332 25248
rect 3384 25236 3390 25288
rect 4617 25279 4675 25285
rect 4617 25245 4629 25279
rect 4663 25276 4675 25279
rect 5534 25276 5540 25288
rect 4663 25248 5540 25276
rect 4663 25245 4675 25248
rect 4617 25239 4675 25245
rect 5534 25236 5540 25248
rect 5592 25236 5598 25288
rect 9309 25279 9367 25285
rect 9309 25245 9321 25279
rect 9355 25276 9367 25279
rect 9674 25276 9680 25288
rect 9355 25248 9680 25276
rect 9355 25245 9367 25248
rect 9309 25239 9367 25245
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 9950 25276 9956 25288
rect 9911 25248 9956 25276
rect 9950 25236 9956 25248
rect 10008 25236 10014 25288
rect 12069 25279 12127 25285
rect 12069 25276 12081 25279
rect 11532 25248 12081 25276
rect 2547 25180 3188 25208
rect 2547 25177 2559 25180
rect 2501 25171 2559 25177
rect 3786 25168 3792 25220
rect 3844 25208 3850 25220
rect 5721 25211 5779 25217
rect 5721 25208 5733 25211
rect 3844 25180 5733 25208
rect 3844 25168 3850 25180
rect 5721 25177 5733 25180
rect 5767 25177 5779 25211
rect 5721 25171 5779 25177
rect 5810 25168 5816 25220
rect 5868 25208 5874 25220
rect 6917 25211 6975 25217
rect 6917 25208 6929 25211
rect 5868 25180 5913 25208
rect 6840 25180 6929 25208
rect 5868 25168 5874 25180
rect 3142 25140 3148 25152
rect 3103 25112 3148 25140
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 4430 25100 4436 25152
rect 4488 25140 4494 25152
rect 4982 25140 4988 25152
rect 4488 25112 4988 25140
rect 4488 25100 4494 25112
rect 4982 25100 4988 25112
rect 5040 25100 5046 25152
rect 5166 25140 5172 25152
rect 5127 25112 5172 25140
rect 5166 25100 5172 25112
rect 5224 25100 5230 25152
rect 5442 25100 5448 25152
rect 5500 25140 5506 25152
rect 6840 25140 6868 25180
rect 6917 25177 6929 25180
rect 6963 25177 6975 25211
rect 6917 25171 6975 25177
rect 7006 25168 7012 25220
rect 7064 25208 7070 25220
rect 7561 25211 7619 25217
rect 7064 25180 7109 25208
rect 7064 25168 7070 25180
rect 7561 25177 7573 25211
rect 7607 25208 7619 25211
rect 8202 25208 8208 25220
rect 7607 25180 8208 25208
rect 7607 25177 7619 25180
rect 7561 25171 7619 25177
rect 8202 25168 8208 25180
rect 8260 25168 8266 25220
rect 8573 25211 8631 25217
rect 8573 25177 8585 25211
rect 8619 25208 8631 25211
rect 9490 25208 9496 25220
rect 8619 25180 9496 25208
rect 8619 25177 8631 25180
rect 8573 25171 8631 25177
rect 9490 25168 9496 25180
rect 9548 25168 9554 25220
rect 11238 25208 11244 25220
rect 11199 25180 11244 25208
rect 11238 25168 11244 25180
rect 11296 25168 11302 25220
rect 8846 25140 8852 25152
rect 5500 25112 8852 25140
rect 5500 25100 5506 25112
rect 8846 25100 8852 25112
rect 8904 25100 8910 25152
rect 9858 25140 9864 25152
rect 9819 25112 9864 25140
rect 9858 25100 9864 25112
rect 9916 25100 9922 25152
rect 10594 25100 10600 25152
rect 10652 25140 10658 25152
rect 11532 25140 11560 25248
rect 12069 25245 12081 25248
rect 12115 25245 12127 25279
rect 13541 25279 13599 25285
rect 13541 25276 13553 25279
rect 12069 25239 12127 25245
rect 12406 25248 13553 25276
rect 11606 25168 11612 25220
rect 11664 25208 11670 25220
rect 11664 25180 12204 25208
rect 11664 25168 11670 25180
rect 10652 25112 11560 25140
rect 12176 25140 12204 25180
rect 12250 25168 12256 25220
rect 12308 25208 12314 25220
rect 12406 25208 12434 25248
rect 13541 25245 13553 25248
rect 13587 25245 13599 25279
rect 13541 25239 13599 25245
rect 13630 25236 13636 25288
rect 13688 25276 13694 25288
rect 13688 25248 13733 25276
rect 13688 25236 13694 25248
rect 14826 25236 14832 25288
rect 14884 25276 14890 25288
rect 15197 25279 15255 25285
rect 15197 25276 15209 25279
rect 14884 25248 15209 25276
rect 14884 25236 14890 25248
rect 15197 25245 15209 25248
rect 15243 25245 15255 25279
rect 15197 25239 15255 25245
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25276 15991 25279
rect 16482 25276 16488 25288
rect 15979 25248 16488 25276
rect 15979 25245 15991 25248
rect 15933 25239 15991 25245
rect 16482 25236 16488 25248
rect 16540 25236 16546 25288
rect 16945 25279 17003 25285
rect 16945 25245 16957 25279
rect 16991 25245 17003 25279
rect 16945 25239 17003 25245
rect 12308 25180 12434 25208
rect 12713 25211 12771 25217
rect 12308 25168 12314 25180
rect 12713 25177 12725 25211
rect 12759 25208 12771 25211
rect 14090 25208 14096 25220
rect 12759 25180 14096 25208
rect 12759 25177 12771 25180
rect 12713 25171 12771 25177
rect 14090 25168 14096 25180
rect 14148 25168 14154 25220
rect 14458 25208 14464 25220
rect 14419 25180 14464 25208
rect 14458 25168 14464 25180
rect 14516 25168 14522 25220
rect 15470 25208 15476 25220
rect 14568 25180 15476 25208
rect 14568 25140 14596 25180
rect 15470 25168 15476 25180
rect 15528 25168 15534 25220
rect 15286 25140 15292 25152
rect 12176 25112 14596 25140
rect 15247 25112 15292 25140
rect 10652 25100 10658 25112
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 16022 25140 16028 25152
rect 15983 25112 16028 25140
rect 16022 25100 16028 25112
rect 16080 25100 16086 25152
rect 16960 25140 16988 25239
rect 17770 25168 17776 25220
rect 17828 25208 17834 25220
rect 20806 25208 20812 25220
rect 17828 25180 17873 25208
rect 17972 25180 19288 25208
rect 20767 25180 20812 25208
rect 17828 25168 17834 25180
rect 17972 25140 18000 25180
rect 19260 25152 19288 25180
rect 20806 25168 20812 25180
rect 20864 25168 20870 25220
rect 16960 25112 18000 25140
rect 18046 25100 18052 25152
rect 18104 25140 18110 25152
rect 18782 25140 18788 25152
rect 18104 25112 18788 25140
rect 18104 25100 18110 25112
rect 18782 25100 18788 25112
rect 18840 25100 18846 25152
rect 19242 25100 19248 25152
rect 19300 25140 19306 25152
rect 19429 25143 19487 25149
rect 19429 25140 19441 25143
rect 19300 25112 19441 25140
rect 19300 25100 19306 25112
rect 19429 25109 19441 25112
rect 19475 25109 19487 25143
rect 19429 25103 19487 25109
rect 1104 25050 36892 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 36892 25050
rect 1104 24976 36892 24998
rect 8128 24908 10640 24936
rect 2133 24871 2191 24877
rect 2133 24837 2145 24871
rect 2179 24868 2191 24871
rect 2222 24868 2228 24880
rect 2179 24840 2228 24868
rect 2179 24837 2191 24840
rect 2133 24831 2191 24837
rect 2222 24828 2228 24840
rect 2280 24828 2286 24880
rect 3786 24868 3792 24880
rect 2700 24840 3792 24868
rect 1946 24692 1952 24744
rect 2004 24732 2010 24744
rect 2225 24735 2283 24741
rect 2225 24732 2237 24735
rect 2004 24704 2237 24732
rect 2004 24692 2010 24704
rect 2225 24701 2237 24704
rect 2271 24732 2283 24735
rect 2700 24732 2728 24840
rect 3786 24828 3792 24840
rect 3844 24828 3850 24880
rect 3878 24828 3884 24880
rect 3936 24868 3942 24880
rect 3936 24840 3981 24868
rect 3936 24828 3942 24840
rect 5534 24828 5540 24880
rect 5592 24868 5598 24880
rect 6638 24868 6644 24880
rect 5592 24840 6644 24868
rect 5592 24828 5598 24840
rect 6638 24828 6644 24840
rect 6696 24828 6702 24880
rect 7282 24828 7288 24880
rect 7340 24868 7346 24880
rect 7926 24868 7932 24880
rect 7340 24840 7932 24868
rect 7340 24828 7346 24840
rect 7926 24828 7932 24840
rect 7984 24868 7990 24880
rect 8128 24868 8156 24908
rect 10502 24868 10508 24880
rect 7984 24840 8156 24868
rect 8588 24840 8892 24868
rect 10463 24840 10508 24868
rect 7984 24828 7990 24840
rect 2774 24760 2780 24812
rect 2832 24800 2838 24812
rect 2832 24772 2877 24800
rect 2832 24760 2838 24772
rect 5626 24760 5632 24812
rect 5684 24800 5690 24812
rect 5813 24803 5871 24809
rect 5813 24800 5825 24803
rect 5684 24772 5825 24800
rect 5684 24760 5690 24772
rect 5813 24769 5825 24772
rect 5859 24769 5871 24803
rect 5813 24763 5871 24769
rect 5902 24760 5908 24812
rect 5960 24800 5966 24812
rect 6549 24803 6607 24809
rect 5960 24772 6005 24800
rect 5960 24760 5966 24772
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 7374 24800 7380 24812
rect 7335 24772 7380 24800
rect 6549 24763 6607 24769
rect 2271 24704 2728 24732
rect 3697 24735 3755 24741
rect 2271 24701 2283 24704
rect 2225 24695 2283 24701
rect 3697 24701 3709 24735
rect 3743 24701 3755 24735
rect 3697 24695 3755 24701
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24732 4031 24735
rect 4019 24704 4660 24732
rect 4019 24701 4031 24704
rect 3973 24695 4031 24701
rect 1673 24667 1731 24673
rect 1673 24633 1685 24667
rect 1719 24664 1731 24667
rect 3712 24664 3740 24695
rect 4522 24664 4528 24676
rect 1719 24636 2774 24664
rect 3712 24636 4528 24664
rect 1719 24633 1731 24636
rect 1673 24627 1731 24633
rect 2746 24596 2774 24636
rect 4522 24624 4528 24636
rect 4580 24624 4586 24676
rect 4430 24596 4436 24608
rect 2746 24568 4436 24596
rect 4430 24556 4436 24568
rect 4488 24556 4494 24608
rect 4632 24605 4660 24704
rect 4982 24692 4988 24744
rect 5040 24732 5046 24744
rect 6564 24732 6592 24763
rect 7374 24760 7380 24772
rect 7432 24760 7438 24812
rect 8036 24809 8064 24840
rect 8021 24803 8079 24809
rect 8021 24769 8033 24803
rect 8067 24769 8079 24803
rect 8021 24763 8079 24769
rect 8110 24760 8116 24812
rect 8168 24800 8174 24812
rect 8588 24800 8616 24840
rect 8168 24772 8616 24800
rect 8168 24760 8174 24772
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 8864 24800 8892 24840
rect 10502 24828 10508 24840
rect 10560 24828 10566 24880
rect 10612 24868 10640 24908
rect 10962 24896 10968 24948
rect 11020 24936 11026 24948
rect 15378 24936 15384 24948
rect 11020 24908 15384 24936
rect 11020 24896 11026 24908
rect 15378 24896 15384 24908
rect 15436 24896 15442 24948
rect 16022 24896 16028 24948
rect 16080 24936 16086 24948
rect 33778 24936 33784 24948
rect 16080 24908 33784 24936
rect 16080 24896 16086 24908
rect 33778 24896 33784 24908
rect 33836 24896 33842 24948
rect 11606 24868 11612 24880
rect 10612 24840 11612 24868
rect 11606 24828 11612 24840
rect 11664 24828 11670 24880
rect 11882 24868 11888 24880
rect 11843 24840 11888 24868
rect 11882 24828 11888 24840
rect 11940 24828 11946 24880
rect 13538 24828 13544 24880
rect 13596 24868 13602 24880
rect 13633 24871 13691 24877
rect 13633 24868 13645 24871
rect 13596 24840 13645 24868
rect 13596 24828 13602 24840
rect 13633 24837 13645 24840
rect 13679 24837 13691 24871
rect 14826 24868 14832 24880
rect 14787 24840 14832 24868
rect 13633 24831 13691 24837
rect 14826 24828 14832 24840
rect 14884 24828 14890 24880
rect 17034 24868 17040 24880
rect 16995 24840 17040 24868
rect 17034 24828 17040 24840
rect 17092 24828 17098 24880
rect 17126 24828 17132 24880
rect 17184 24868 17190 24880
rect 17770 24868 17776 24880
rect 17184 24840 17776 24868
rect 17184 24828 17190 24840
rect 17770 24828 17776 24840
rect 17828 24828 17834 24880
rect 9401 24803 9459 24809
rect 9401 24800 9413 24803
rect 8720 24772 8765 24800
rect 8864 24772 9413 24800
rect 8720 24760 8726 24772
rect 9401 24769 9413 24772
rect 9447 24769 9459 24803
rect 9401 24763 9459 24769
rect 9493 24803 9551 24809
rect 9493 24769 9505 24803
rect 9539 24800 9551 24803
rect 9950 24800 9956 24812
rect 9539 24772 9956 24800
rect 9539 24769 9551 24772
rect 9493 24763 9551 24769
rect 9950 24760 9956 24772
rect 10008 24760 10014 24812
rect 14182 24760 14188 24812
rect 14240 24800 14246 24812
rect 18506 24800 18512 24812
rect 14240 24772 14285 24800
rect 18467 24772 18512 24800
rect 14240 24760 14246 24772
rect 18506 24760 18512 24772
rect 18564 24760 18570 24812
rect 18598 24760 18604 24812
rect 18656 24800 18662 24812
rect 18656 24772 18701 24800
rect 18656 24760 18662 24772
rect 18782 24760 18788 24812
rect 18840 24800 18846 24812
rect 21082 24800 21088 24812
rect 18840 24772 21088 24800
rect 18840 24760 18846 24772
rect 21082 24760 21088 24772
rect 21140 24760 21146 24812
rect 5040 24704 6592 24732
rect 6641 24735 6699 24741
rect 5040 24692 5046 24704
rect 6641 24701 6653 24735
rect 6687 24732 6699 24735
rect 6730 24732 6736 24744
rect 6687 24704 6736 24732
rect 6687 24701 6699 24704
rect 6641 24695 6699 24701
rect 6730 24692 6736 24704
rect 6788 24692 6794 24744
rect 7469 24735 7527 24741
rect 7469 24701 7481 24735
rect 7515 24732 7527 24735
rect 7515 24704 10548 24732
rect 7515 24701 7527 24704
rect 7469 24695 7527 24701
rect 5353 24667 5411 24673
rect 5353 24633 5365 24667
rect 5399 24664 5411 24667
rect 6178 24664 6184 24676
rect 5399 24636 6184 24664
rect 5399 24633 5411 24636
rect 5353 24627 5411 24633
rect 6178 24624 6184 24636
rect 6236 24624 6242 24676
rect 6362 24624 6368 24676
rect 6420 24664 6426 24676
rect 8662 24664 8668 24676
rect 6420 24636 8668 24664
rect 6420 24624 6426 24636
rect 8662 24624 8668 24636
rect 8720 24624 8726 24676
rect 8757 24667 8815 24673
rect 8757 24633 8769 24667
rect 8803 24664 8815 24667
rect 8803 24636 9996 24664
rect 8803 24633 8815 24636
rect 8757 24627 8815 24633
rect 4617 24599 4675 24605
rect 4617 24565 4629 24599
rect 4663 24596 4675 24599
rect 4798 24596 4804 24608
rect 4663 24568 4804 24596
rect 4663 24565 4675 24568
rect 4617 24559 4675 24565
rect 4798 24556 4804 24568
rect 4856 24556 4862 24608
rect 4890 24556 4896 24608
rect 4948 24596 4954 24608
rect 8018 24596 8024 24608
rect 4948 24568 8024 24596
rect 4948 24556 4954 24568
rect 8018 24556 8024 24568
rect 8076 24556 8082 24608
rect 8113 24599 8171 24605
rect 8113 24565 8125 24599
rect 8159 24596 8171 24599
rect 8938 24596 8944 24608
rect 8159 24568 8944 24596
rect 8159 24565 8171 24568
rect 8113 24559 8171 24565
rect 8938 24556 8944 24568
rect 8996 24556 9002 24608
rect 9968 24596 9996 24636
rect 10042 24624 10048 24676
rect 10100 24664 10106 24676
rect 10520 24664 10548 24704
rect 10594 24692 10600 24744
rect 10652 24732 10658 24744
rect 10652 24704 10697 24732
rect 10652 24692 10658 24704
rect 11330 24692 11336 24744
rect 11388 24732 11394 24744
rect 11793 24735 11851 24741
rect 11793 24732 11805 24735
rect 11388 24704 11805 24732
rect 11388 24692 11394 24704
rect 11793 24701 11805 24704
rect 11839 24701 11851 24735
rect 13262 24732 13268 24744
rect 11793 24695 11851 24701
rect 11900 24704 13268 24732
rect 11900 24664 11928 24704
rect 13262 24692 13268 24704
rect 13320 24692 13326 24744
rect 13354 24692 13360 24744
rect 13412 24732 13418 24744
rect 13541 24735 13599 24741
rect 13541 24732 13553 24735
rect 13412 24704 13553 24732
rect 13412 24692 13418 24704
rect 13541 24701 13553 24704
rect 13587 24701 13599 24735
rect 14734 24732 14740 24744
rect 14695 24704 14740 24732
rect 13541 24695 13599 24701
rect 14734 24692 14740 24704
rect 14792 24692 14798 24744
rect 15749 24735 15807 24741
rect 15749 24701 15761 24735
rect 15795 24732 15807 24735
rect 16945 24735 17003 24741
rect 15795 24704 16574 24732
rect 15795 24701 15807 24704
rect 15749 24695 15807 24701
rect 12342 24664 12348 24676
rect 10100 24636 10145 24664
rect 10520 24636 11928 24664
rect 12303 24636 12348 24664
rect 10100 24624 10106 24636
rect 12342 24624 12348 24636
rect 12400 24624 12406 24676
rect 14458 24664 14464 24676
rect 12820 24636 14464 24664
rect 12820 24596 12848 24636
rect 14458 24624 14464 24636
rect 14516 24624 14522 24676
rect 16546 24664 16574 24704
rect 16945 24701 16957 24735
rect 16991 24732 17003 24735
rect 17126 24732 17132 24744
rect 16991 24704 17132 24732
rect 16991 24701 17003 24704
rect 16945 24695 17003 24701
rect 17126 24692 17132 24704
rect 17184 24692 17190 24744
rect 17221 24735 17279 24741
rect 17221 24701 17233 24735
rect 17267 24732 17279 24735
rect 17310 24732 17316 24744
rect 17267 24704 17316 24732
rect 17267 24701 17279 24704
rect 17221 24695 17279 24701
rect 17236 24664 17264 24695
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 18616 24732 18644 24760
rect 19061 24735 19119 24741
rect 19061 24732 19073 24735
rect 18616 24704 19073 24732
rect 19061 24701 19073 24704
rect 19107 24701 19119 24735
rect 19061 24695 19119 24701
rect 35894 24692 35900 24744
rect 35952 24732 35958 24744
rect 36081 24735 36139 24741
rect 36081 24732 36093 24735
rect 35952 24704 36093 24732
rect 35952 24692 35958 24704
rect 36081 24701 36093 24704
rect 36127 24701 36139 24735
rect 36354 24732 36360 24744
rect 36315 24704 36360 24732
rect 36081 24695 36139 24701
rect 36354 24692 36360 24704
rect 36412 24692 36418 24744
rect 16546 24636 17264 24664
rect 12986 24596 12992 24608
rect 9968 24568 12848 24596
rect 12947 24568 12992 24596
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 16301 24599 16359 24605
rect 16301 24565 16313 24599
rect 16347 24596 16359 24599
rect 17310 24596 17316 24608
rect 16347 24568 17316 24596
rect 16347 24565 16359 24568
rect 16301 24559 16359 24565
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 19242 24556 19248 24608
rect 19300 24596 19306 24608
rect 19705 24599 19763 24605
rect 19705 24596 19717 24599
rect 19300 24568 19717 24596
rect 19300 24556 19306 24568
rect 19705 24565 19717 24568
rect 19751 24565 19763 24599
rect 19705 24559 19763 24565
rect 1104 24506 36892 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 36892 24506
rect 1104 24432 36892 24454
rect 2130 24352 2136 24404
rect 2188 24392 2194 24404
rect 2225 24395 2283 24401
rect 2225 24392 2237 24395
rect 2188 24364 2237 24392
rect 2188 24352 2194 24364
rect 2225 24361 2237 24364
rect 2271 24361 2283 24395
rect 2225 24355 2283 24361
rect 3326 24352 3332 24404
rect 3384 24392 3390 24404
rect 3973 24395 4031 24401
rect 3973 24392 3985 24395
rect 3384 24364 3985 24392
rect 3384 24352 3390 24364
rect 3973 24361 3985 24364
rect 4019 24361 4031 24395
rect 3973 24355 4031 24361
rect 5810 24352 5816 24404
rect 5868 24392 5874 24404
rect 6365 24395 6423 24401
rect 6365 24392 6377 24395
rect 5868 24364 6377 24392
rect 5868 24352 5874 24364
rect 6365 24361 6377 24364
rect 6411 24361 6423 24395
rect 7006 24392 7012 24404
rect 6967 24364 7012 24392
rect 6365 24355 6423 24361
rect 7006 24352 7012 24364
rect 7064 24352 7070 24404
rect 7098 24352 7104 24404
rect 7156 24392 7162 24404
rect 13538 24392 13544 24404
rect 7156 24364 8524 24392
rect 7156 24352 7162 24364
rect 1394 24284 1400 24336
rect 1452 24324 1458 24336
rect 8496 24324 8524 24364
rect 9324 24364 13544 24392
rect 9214 24324 9220 24336
rect 1452 24296 8432 24324
rect 8496 24296 9220 24324
rect 1452 24284 1458 24296
rect 1762 24216 1768 24268
rect 1820 24256 1826 24268
rect 2869 24259 2927 24265
rect 1820 24228 2820 24256
rect 1820 24216 1826 24228
rect 1946 24148 1952 24200
rect 2004 24188 2010 24200
rect 2792 24197 2820 24228
rect 2869 24225 2881 24259
rect 2915 24256 2927 24259
rect 4890 24256 4896 24268
rect 2915 24228 4896 24256
rect 2915 24225 2927 24228
rect 2869 24219 2927 24225
rect 4890 24216 4896 24228
rect 4948 24216 4954 24268
rect 5258 24216 5264 24268
rect 5316 24256 5322 24268
rect 5316 24228 7788 24256
rect 5316 24216 5322 24228
rect 2317 24191 2375 24197
rect 2317 24188 2329 24191
rect 2004 24160 2329 24188
rect 2004 24148 2010 24160
rect 2317 24157 2329 24160
rect 2363 24157 2375 24191
rect 2317 24151 2375 24157
rect 2777 24191 2835 24197
rect 2777 24157 2789 24191
rect 2823 24188 2835 24191
rect 4157 24191 4215 24197
rect 4157 24188 4169 24191
rect 2823 24160 4169 24188
rect 2823 24157 2835 24160
rect 2777 24151 2835 24157
rect 4157 24157 4169 24160
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 5074 24148 5080 24200
rect 5132 24188 5138 24200
rect 5169 24191 5227 24197
rect 5169 24188 5181 24191
rect 5132 24160 5181 24188
rect 5132 24148 5138 24160
rect 5169 24157 5181 24160
rect 5215 24157 5227 24191
rect 5169 24151 5227 24157
rect 6457 24191 6515 24197
rect 6457 24157 6469 24191
rect 6503 24188 6515 24191
rect 6730 24188 6736 24200
rect 6503 24160 6736 24188
rect 6503 24157 6515 24160
rect 6457 24151 6515 24157
rect 6730 24148 6736 24160
rect 6788 24148 6794 24200
rect 7098 24188 7104 24200
rect 7059 24160 7104 24188
rect 7098 24148 7104 24160
rect 7156 24148 7162 24200
rect 7760 24197 7788 24228
rect 7745 24191 7803 24197
rect 7745 24157 7757 24191
rect 7791 24157 7803 24191
rect 7745 24151 7803 24157
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 8404 24197 8432 24296
rect 9214 24284 9220 24296
rect 9272 24284 9278 24336
rect 8481 24259 8539 24265
rect 8481 24225 8493 24259
rect 8527 24256 8539 24259
rect 9324 24256 9352 24364
rect 13538 24352 13544 24364
rect 13596 24352 13602 24404
rect 15562 24392 15568 24404
rect 13740 24364 15568 24392
rect 13740 24336 13768 24364
rect 15562 24352 15568 24364
rect 15620 24352 15626 24404
rect 20806 24352 20812 24404
rect 20864 24392 20870 24404
rect 20901 24395 20959 24401
rect 20901 24392 20913 24395
rect 20864 24364 20913 24392
rect 20864 24352 20870 24364
rect 20901 24361 20913 24364
rect 20947 24361 20959 24395
rect 36354 24392 36360 24404
rect 36315 24364 36360 24392
rect 20901 24355 20959 24361
rect 36354 24352 36360 24364
rect 36412 24352 36418 24404
rect 10045 24327 10103 24333
rect 10045 24293 10057 24327
rect 10091 24324 10103 24327
rect 12710 24324 12716 24336
rect 10091 24296 12716 24324
rect 10091 24293 10103 24296
rect 10045 24287 10103 24293
rect 12710 24284 12716 24296
rect 12768 24284 12774 24336
rect 12986 24284 12992 24336
rect 13044 24324 13050 24336
rect 13722 24324 13728 24336
rect 13044 24296 13728 24324
rect 13044 24284 13050 24296
rect 13722 24284 13728 24296
rect 13780 24284 13786 24336
rect 14734 24284 14740 24336
rect 14792 24324 14798 24336
rect 14792 24296 18276 24324
rect 14792 24284 14798 24296
rect 9490 24256 9496 24268
rect 8527 24228 9352 24256
rect 9451 24228 9496 24256
rect 8527 24225 8539 24228
rect 8481 24219 8539 24225
rect 9490 24216 9496 24228
rect 9548 24216 9554 24268
rect 10689 24259 10747 24265
rect 10689 24225 10701 24259
rect 10735 24256 10747 24259
rect 11054 24256 11060 24268
rect 10735 24228 11060 24256
rect 10735 24225 10747 24228
rect 10689 24219 10747 24225
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 11333 24259 11391 24265
rect 11333 24225 11345 24259
rect 11379 24256 11391 24259
rect 12158 24256 12164 24268
rect 11379 24228 12164 24256
rect 11379 24225 11391 24228
rect 11333 24219 11391 24225
rect 12158 24216 12164 24228
rect 12216 24216 12222 24268
rect 12434 24256 12440 24268
rect 12395 24228 12440 24256
rect 12434 24216 12440 24228
rect 12492 24256 12498 24268
rect 12802 24256 12808 24268
rect 12492 24228 12808 24256
rect 12492 24216 12498 24228
rect 12802 24216 12808 24228
rect 12860 24256 12866 24268
rect 13081 24259 13139 24265
rect 13081 24256 13093 24259
rect 12860 24228 13093 24256
rect 12860 24216 12866 24228
rect 13081 24225 13093 24228
rect 13127 24225 13139 24259
rect 13081 24219 13139 24225
rect 13170 24216 13176 24268
rect 13228 24256 13234 24268
rect 13357 24259 13415 24265
rect 13357 24256 13369 24259
rect 13228 24228 13369 24256
rect 13228 24216 13234 24228
rect 13357 24225 13369 24228
rect 13403 24225 13415 24259
rect 13357 24219 13415 24225
rect 14182 24216 14188 24268
rect 14240 24256 14246 24268
rect 14645 24259 14703 24265
rect 14645 24256 14657 24259
rect 14240 24228 14657 24256
rect 14240 24216 14246 24228
rect 14645 24225 14657 24228
rect 14691 24225 14703 24259
rect 14645 24219 14703 24225
rect 15565 24259 15623 24265
rect 15565 24225 15577 24259
rect 15611 24256 15623 24259
rect 16482 24256 16488 24268
rect 15611 24228 16488 24256
rect 15611 24225 15623 24228
rect 15565 24219 15623 24225
rect 16482 24216 16488 24228
rect 16540 24216 16546 24268
rect 16669 24259 16727 24265
rect 16669 24225 16681 24259
rect 16715 24256 16727 24259
rect 17494 24256 17500 24268
rect 16715 24228 17500 24256
rect 16715 24225 16727 24228
rect 16669 24219 16727 24225
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 17957 24259 18015 24265
rect 17957 24225 17969 24259
rect 18003 24256 18015 24259
rect 18138 24256 18144 24268
rect 18003 24228 18144 24256
rect 18003 24225 18015 24228
rect 17957 24219 18015 24225
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 18248 24265 18276 24296
rect 18233 24259 18291 24265
rect 18233 24225 18245 24259
rect 18279 24225 18291 24259
rect 18233 24219 18291 24225
rect 8389 24191 8447 24197
rect 7892 24160 7937 24188
rect 7892 24148 7898 24160
rect 8389 24157 8401 24191
rect 8435 24157 8447 24191
rect 8389 24151 8447 24157
rect 17218 24148 17224 24200
rect 17276 24188 17282 24200
rect 17405 24191 17463 24197
rect 17405 24188 17417 24191
rect 17276 24160 17417 24188
rect 17276 24148 17282 24160
rect 17405 24157 17417 24160
rect 17451 24157 17463 24191
rect 17405 24151 17463 24157
rect 5261 24123 5319 24129
rect 5261 24089 5273 24123
rect 5307 24120 5319 24123
rect 9585 24123 9643 24129
rect 5307 24092 9352 24120
rect 5307 24089 5319 24092
rect 5261 24083 5319 24089
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 4614 24052 4620 24064
rect 4575 24024 4620 24052
rect 4614 24012 4620 24024
rect 4672 24012 4678 24064
rect 5350 24012 5356 24064
rect 5408 24052 5414 24064
rect 8478 24052 8484 24064
rect 5408 24024 8484 24052
rect 5408 24012 5414 24024
rect 8478 24012 8484 24024
rect 8536 24012 8542 24064
rect 9324 24052 9352 24092
rect 9585 24089 9597 24123
rect 9631 24089 9643 24123
rect 9585 24083 9643 24089
rect 9600 24052 9628 24083
rect 10778 24080 10784 24132
rect 10836 24120 10842 24132
rect 12345 24123 12403 24129
rect 10836 24092 10881 24120
rect 10836 24080 10842 24092
rect 12345 24089 12357 24123
rect 12391 24089 12403 24123
rect 12345 24083 12403 24089
rect 13173 24123 13231 24129
rect 13173 24089 13185 24123
rect 13219 24089 13231 24123
rect 13173 24083 13231 24089
rect 9324 24024 9628 24052
rect 10042 24012 10048 24064
rect 10100 24052 10106 24064
rect 10870 24052 10876 24064
rect 10100 24024 10876 24052
rect 10100 24012 10106 24024
rect 10870 24012 10876 24024
rect 10928 24012 10934 24064
rect 12360 24052 12388 24083
rect 12618 24052 12624 24064
rect 12360 24024 12624 24052
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 13188 24052 13216 24083
rect 14090 24080 14096 24132
rect 14148 24120 14154 24132
rect 14369 24123 14427 24129
rect 14369 24120 14381 24123
rect 14148 24092 14381 24120
rect 14148 24080 14154 24092
rect 14369 24089 14381 24092
rect 14415 24089 14427 24123
rect 14369 24083 14427 24089
rect 14458 24080 14464 24132
rect 14516 24120 14522 24132
rect 14516 24092 14561 24120
rect 14516 24080 14522 24092
rect 15930 24080 15936 24132
rect 15988 24120 15994 24132
rect 16025 24123 16083 24129
rect 16025 24120 16037 24123
rect 15988 24092 16037 24120
rect 15988 24080 15994 24092
rect 16025 24089 16037 24092
rect 16071 24089 16083 24123
rect 16025 24083 16083 24089
rect 16574 24080 16580 24132
rect 16632 24120 16638 24132
rect 17420 24120 17448 24151
rect 18782 24148 18788 24200
rect 18840 24188 18846 24200
rect 19242 24188 19248 24200
rect 18840 24160 19248 24188
rect 18840 24148 18846 24160
rect 19242 24148 19248 24160
rect 19300 24188 19306 24200
rect 19889 24191 19947 24197
rect 19889 24188 19901 24191
rect 19300 24160 19901 24188
rect 19300 24148 19306 24160
rect 19889 24157 19901 24160
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 20993 24191 21051 24197
rect 20993 24157 21005 24191
rect 21039 24188 21051 24191
rect 21039 24160 21128 24188
rect 21039 24157 21051 24160
rect 20993 24151 21051 24157
rect 17954 24120 17960 24132
rect 16632 24092 16677 24120
rect 17420 24092 17960 24120
rect 16632 24080 16638 24092
rect 17954 24080 17960 24092
rect 18012 24080 18018 24132
rect 18046 24080 18052 24132
rect 18104 24120 18110 24132
rect 18104 24092 18149 24120
rect 18104 24080 18110 24092
rect 21100 24064 21128 24160
rect 24670 24080 24676 24132
rect 24728 24120 24734 24132
rect 34790 24120 34796 24132
rect 24728 24092 34796 24120
rect 24728 24080 24734 24092
rect 34790 24080 34796 24092
rect 34848 24080 34854 24132
rect 13814 24052 13820 24064
rect 13188 24024 13820 24052
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 16114 24012 16120 24064
rect 16172 24052 16178 24064
rect 17313 24055 17371 24061
rect 17313 24052 17325 24055
rect 16172 24024 17325 24052
rect 16172 24012 16178 24024
rect 17313 24021 17325 24024
rect 17359 24021 17371 24055
rect 17313 24015 17371 24021
rect 19981 24055 20039 24061
rect 19981 24021 19993 24055
rect 20027 24052 20039 24055
rect 20254 24052 20260 24064
rect 20027 24024 20260 24052
rect 20027 24021 20039 24024
rect 19981 24015 20039 24021
rect 20254 24012 20260 24024
rect 20312 24012 20318 24064
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 21453 24055 21511 24061
rect 21453 24052 21465 24055
rect 21140 24024 21465 24052
rect 21140 24012 21146 24024
rect 21453 24021 21465 24024
rect 21499 24021 21511 24055
rect 21453 24015 21511 24021
rect 1104 23962 36892 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 36892 23962
rect 1104 23888 36892 23910
rect 2222 23808 2228 23860
rect 2280 23848 2286 23860
rect 3234 23848 3240 23860
rect 2280 23820 3240 23848
rect 2280 23808 2286 23820
rect 3234 23808 3240 23820
rect 3292 23808 3298 23860
rect 5810 23848 5816 23860
rect 3344 23820 5816 23848
rect 3344 23780 3372 23820
rect 5810 23808 5816 23820
rect 5868 23808 5874 23860
rect 6454 23808 6460 23860
rect 6512 23848 6518 23860
rect 7098 23848 7104 23860
rect 6512 23820 7104 23848
rect 6512 23808 6518 23820
rect 7098 23808 7104 23820
rect 7156 23808 7162 23860
rect 10042 23848 10048 23860
rect 8220 23820 10048 23848
rect 5445 23783 5503 23789
rect 5445 23780 5457 23783
rect 2240 23752 3372 23780
rect 3436 23752 5457 23780
rect 2240 23721 2268 23752
rect 2225 23715 2283 23721
rect 2225 23681 2237 23715
rect 2271 23681 2283 23715
rect 2225 23675 2283 23681
rect 2685 23715 2743 23721
rect 2685 23681 2697 23715
rect 2731 23681 2743 23715
rect 2685 23675 2743 23681
rect 2777 23715 2835 23721
rect 2777 23681 2789 23715
rect 2823 23712 2835 23715
rect 3436 23712 3464 23752
rect 5445 23749 5457 23752
rect 5491 23749 5503 23783
rect 5445 23743 5503 23749
rect 6822 23740 6828 23792
rect 6880 23780 6886 23792
rect 8220 23789 8248 23820
rect 10042 23808 10048 23820
rect 10100 23808 10106 23860
rect 11790 23848 11796 23860
rect 10152 23820 11796 23848
rect 8113 23783 8171 23789
rect 8113 23780 8125 23783
rect 6880 23752 8125 23780
rect 6880 23740 6886 23752
rect 8113 23749 8125 23752
rect 8159 23749 8171 23783
rect 8113 23743 8171 23749
rect 8205 23783 8263 23789
rect 8205 23749 8217 23783
rect 8251 23749 8263 23783
rect 8938 23780 8944 23792
rect 8899 23752 8944 23780
rect 8205 23743 8263 23749
rect 8938 23740 8944 23752
rect 8996 23740 9002 23792
rect 9490 23780 9496 23792
rect 9403 23752 9496 23780
rect 9490 23740 9496 23752
rect 9548 23780 9554 23792
rect 10152 23780 10180 23820
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 13814 23848 13820 23860
rect 12728 23820 13820 23848
rect 10962 23780 10968 23792
rect 9548 23752 10180 23780
rect 10923 23752 10968 23780
rect 9548 23740 9554 23752
rect 10962 23740 10968 23752
rect 11020 23740 11026 23792
rect 11054 23740 11060 23792
rect 11112 23780 11118 23792
rect 12728 23789 12756 23820
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 14001 23851 14059 23857
rect 14001 23817 14013 23851
rect 14047 23848 14059 23851
rect 14090 23848 14096 23860
rect 14047 23820 14096 23848
rect 14047 23817 14059 23820
rect 14001 23811 14059 23817
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 27798 23848 27804 23860
rect 27759 23820 27804 23848
rect 27798 23808 27804 23820
rect 27856 23808 27862 23860
rect 12713 23783 12771 23789
rect 11112 23752 11157 23780
rect 11112 23740 11118 23752
rect 12713 23749 12725 23783
rect 12759 23749 12771 23783
rect 12713 23743 12771 23749
rect 12802 23740 12808 23792
rect 12860 23780 12866 23792
rect 15930 23780 15936 23792
rect 12860 23752 12905 23780
rect 13004 23752 15936 23780
rect 12860 23740 12866 23752
rect 2823 23684 3464 23712
rect 3513 23715 3571 23721
rect 2823 23681 2835 23684
rect 2777 23675 2835 23681
rect 3513 23681 3525 23715
rect 3559 23712 3571 23715
rect 3786 23712 3792 23724
rect 3559 23684 3792 23712
rect 3559 23681 3571 23684
rect 3513 23675 3571 23681
rect 2038 23604 2044 23656
rect 2096 23644 2102 23656
rect 2700 23644 2728 23675
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 3973 23715 4031 23721
rect 3973 23710 3985 23715
rect 3896 23682 3985 23710
rect 3896 23644 3924 23682
rect 3973 23681 3985 23682
rect 4019 23681 4031 23715
rect 3973 23675 4031 23681
rect 6917 23715 6975 23721
rect 6917 23681 6929 23715
rect 6963 23712 6975 23715
rect 7006 23712 7012 23724
rect 6963 23684 7012 23712
rect 6963 23681 6975 23684
rect 6917 23675 6975 23681
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 12161 23715 12219 23721
rect 12161 23712 12173 23715
rect 11348 23684 12173 23712
rect 11348 23656 11376 23684
rect 12161 23681 12173 23684
rect 12207 23681 12219 23715
rect 12161 23675 12219 23681
rect 5350 23644 5356 23656
rect 2096 23616 2728 23644
rect 3160 23616 3924 23644
rect 5311 23616 5356 23644
rect 2096 23604 2102 23616
rect 1670 23536 1676 23588
rect 1728 23576 1734 23588
rect 3160 23576 3188 23616
rect 5350 23604 5356 23616
rect 5408 23604 5414 23656
rect 5718 23644 5724 23656
rect 5679 23616 5724 23644
rect 5718 23604 5724 23616
rect 5776 23644 5782 23656
rect 7561 23647 7619 23653
rect 7561 23644 7573 23647
rect 5776 23616 7573 23644
rect 5776 23604 5782 23616
rect 7561 23613 7573 23616
rect 7607 23613 7619 23647
rect 7561 23607 7619 23613
rect 8018 23604 8024 23656
rect 8076 23644 8082 23656
rect 8849 23647 8907 23653
rect 8849 23644 8861 23647
rect 8076 23616 8861 23644
rect 8076 23604 8082 23616
rect 8849 23613 8861 23616
rect 8895 23613 8907 23647
rect 8849 23607 8907 23613
rect 1728 23548 3188 23576
rect 1728 23536 1734 23548
rect 3234 23536 3240 23588
rect 3292 23576 3298 23588
rect 3421 23579 3479 23585
rect 3421 23576 3433 23579
rect 3292 23548 3433 23576
rect 3292 23536 3298 23548
rect 3421 23545 3433 23548
rect 3467 23545 3479 23579
rect 3421 23539 3479 23545
rect 3510 23536 3516 23588
rect 3568 23576 3574 23588
rect 4709 23579 4767 23585
rect 4709 23576 4721 23579
rect 3568 23548 4721 23576
rect 3568 23536 3574 23548
rect 4709 23545 4721 23548
rect 4755 23545 4767 23579
rect 4709 23539 4767 23545
rect 4798 23536 4804 23588
rect 4856 23576 4862 23588
rect 8662 23576 8668 23588
rect 4856 23548 8668 23576
rect 4856 23536 4862 23548
rect 8662 23536 8668 23548
rect 8720 23536 8726 23588
rect 8864 23576 8892 23607
rect 8938 23604 8944 23656
rect 8996 23644 9002 23656
rect 10410 23644 10416 23656
rect 8996 23616 10416 23644
rect 8996 23604 9002 23616
rect 10410 23604 10416 23616
rect 10468 23604 10474 23656
rect 10781 23647 10839 23653
rect 10781 23613 10793 23647
rect 10827 23644 10839 23647
rect 11330 23644 11336 23656
rect 10827 23616 11336 23644
rect 10827 23613 10839 23616
rect 10781 23607 10839 23613
rect 11330 23604 11336 23616
rect 11388 23604 11394 23656
rect 11698 23604 11704 23656
rect 11756 23644 11762 23656
rect 12342 23644 12348 23656
rect 11756 23632 12112 23644
rect 12176 23632 12348 23644
rect 11756 23616 12348 23632
rect 11756 23604 11762 23616
rect 12084 23604 12204 23616
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 13004 23644 13032 23752
rect 15930 23740 15936 23752
rect 15988 23740 15994 23792
rect 16114 23780 16120 23792
rect 16075 23752 16120 23780
rect 16114 23740 16120 23752
rect 16172 23740 16178 23792
rect 17034 23780 17040 23792
rect 16995 23752 17040 23780
rect 17034 23740 17040 23752
rect 17092 23740 17098 23792
rect 17402 23740 17408 23792
rect 17460 23780 17466 23792
rect 17589 23783 17647 23789
rect 17589 23780 17601 23783
rect 17460 23752 17601 23780
rect 17460 23740 17466 23752
rect 17589 23749 17601 23752
rect 17635 23780 17647 23783
rect 19705 23783 19763 23789
rect 19705 23780 19717 23783
rect 17635 23752 19717 23780
rect 17635 23749 17647 23752
rect 17589 23743 17647 23749
rect 19705 23749 19717 23752
rect 19751 23749 19763 23783
rect 20254 23780 20260 23792
rect 20215 23752 20260 23780
rect 19705 23743 19763 23749
rect 20254 23740 20260 23752
rect 20312 23740 20318 23792
rect 13078 23672 13084 23724
rect 13136 23712 13142 23724
rect 13357 23715 13415 23721
rect 13357 23712 13369 23715
rect 13136 23684 13369 23712
rect 13136 23672 13142 23684
rect 13357 23681 13369 23684
rect 13403 23681 13415 23715
rect 13357 23675 13415 23681
rect 18782 23672 18788 23724
rect 18840 23712 18846 23724
rect 19061 23715 19119 23721
rect 19061 23712 19073 23715
rect 18840 23684 19073 23712
rect 18840 23672 18846 23684
rect 19061 23681 19073 23684
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 22189 23715 22247 23721
rect 22189 23681 22201 23715
rect 22235 23712 22247 23715
rect 27614 23712 27620 23724
rect 22235 23684 22784 23712
rect 27575 23684 27620 23712
rect 22235 23681 22247 23684
rect 22189 23675 22247 23681
rect 12492 23616 13032 23644
rect 13449 23647 13507 23653
rect 12492 23604 12498 23616
rect 13449 23613 13461 23647
rect 13495 23644 13507 23647
rect 14461 23647 14519 23653
rect 14461 23644 14473 23647
rect 13495 23616 14473 23644
rect 13495 23613 13507 23616
rect 13449 23607 13507 23613
rect 14461 23613 14473 23616
rect 14507 23613 14519 23647
rect 14461 23607 14519 23613
rect 14645 23647 14703 23653
rect 14645 23613 14657 23647
rect 14691 23644 14703 23647
rect 14918 23644 14924 23656
rect 14691 23616 14924 23644
rect 14691 23613 14703 23616
rect 14645 23607 14703 23613
rect 14918 23604 14924 23616
rect 14976 23604 14982 23656
rect 15933 23647 15991 23653
rect 15933 23613 15945 23647
rect 15979 23613 15991 23647
rect 16206 23644 16212 23656
rect 16167 23616 16212 23644
rect 15933 23607 15991 23613
rect 10502 23576 10508 23588
rect 8864 23548 10508 23576
rect 10502 23536 10508 23548
rect 10560 23536 10566 23588
rect 11790 23536 11796 23588
rect 11848 23576 11854 23588
rect 15948 23576 15976 23607
rect 16206 23604 16212 23616
rect 16264 23604 16270 23656
rect 16945 23647 17003 23653
rect 16945 23613 16957 23647
rect 16991 23644 17003 23647
rect 17218 23644 17224 23656
rect 16991 23616 17224 23644
rect 16991 23613 17003 23616
rect 16945 23607 17003 23613
rect 17218 23604 17224 23616
rect 17276 23644 17282 23656
rect 18601 23647 18659 23653
rect 17276 23616 18552 23644
rect 17276 23604 17282 23616
rect 18524 23576 18552 23616
rect 18601 23613 18613 23647
rect 18647 23644 18659 23647
rect 19518 23644 19524 23656
rect 18647 23616 19524 23644
rect 18647 23613 18659 23616
rect 18601 23607 18659 23613
rect 19518 23604 19524 23616
rect 19576 23604 19582 23656
rect 20349 23647 20407 23653
rect 20349 23613 20361 23647
rect 20395 23644 20407 23647
rect 21266 23644 21272 23656
rect 20395 23616 21272 23644
rect 20395 23613 20407 23616
rect 20349 23607 20407 23613
rect 21266 23604 21272 23616
rect 21324 23604 21330 23656
rect 11848 23548 16574 23576
rect 18524 23548 19748 23576
rect 11848 23536 11854 23548
rect 2133 23511 2191 23517
rect 2133 23477 2145 23511
rect 2179 23508 2191 23511
rect 3878 23508 3884 23520
rect 2179 23480 3884 23508
rect 2179 23477 2191 23480
rect 2133 23471 2191 23477
rect 3878 23468 3884 23480
rect 3936 23468 3942 23520
rect 4065 23511 4123 23517
rect 4065 23477 4077 23511
rect 4111 23508 4123 23511
rect 5442 23508 5448 23520
rect 4111 23480 5448 23508
rect 4111 23477 4123 23480
rect 4065 23471 4123 23477
rect 5442 23468 5448 23480
rect 5500 23468 5506 23520
rect 7009 23511 7067 23517
rect 7009 23477 7021 23511
rect 7055 23508 7067 23511
rect 14826 23508 14832 23520
rect 7055 23480 14832 23508
rect 7055 23477 7067 23480
rect 7009 23471 7067 23477
rect 14826 23468 14832 23480
rect 14884 23468 14890 23520
rect 16546 23508 16574 23548
rect 17494 23508 17500 23520
rect 16546 23480 17500 23508
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 19153 23511 19211 23517
rect 19153 23477 19165 23511
rect 19199 23508 19211 23511
rect 19610 23508 19616 23520
rect 19199 23480 19616 23508
rect 19199 23477 19211 23480
rect 19153 23471 19211 23477
rect 19610 23468 19616 23480
rect 19668 23468 19674 23520
rect 19720 23508 19748 23548
rect 22756 23517 22784 23684
rect 27614 23672 27620 23684
rect 27672 23712 27678 23724
rect 28261 23715 28319 23721
rect 28261 23712 28273 23715
rect 27672 23684 28273 23712
rect 27672 23672 27678 23684
rect 28261 23681 28273 23684
rect 28307 23681 28319 23715
rect 28261 23675 28319 23681
rect 22097 23511 22155 23517
rect 22097 23508 22109 23511
rect 19720 23480 22109 23508
rect 22097 23477 22109 23480
rect 22143 23477 22155 23511
rect 22097 23471 22155 23477
rect 22741 23511 22799 23517
rect 22741 23477 22753 23511
rect 22787 23508 22799 23511
rect 23750 23508 23756 23520
rect 22787 23480 23756 23508
rect 22787 23477 22799 23480
rect 22741 23471 22799 23477
rect 23750 23468 23756 23480
rect 23808 23468 23814 23520
rect 1104 23418 36892 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 36892 23418
rect 1104 23344 36892 23366
rect 2133 23307 2191 23313
rect 2133 23273 2145 23307
rect 2179 23304 2191 23307
rect 2406 23304 2412 23316
rect 2179 23276 2412 23304
rect 2179 23273 2191 23276
rect 2133 23267 2191 23273
rect 2406 23264 2412 23276
rect 2464 23264 2470 23316
rect 3421 23307 3479 23313
rect 3421 23273 3433 23307
rect 3467 23304 3479 23307
rect 3510 23304 3516 23316
rect 3467 23276 3516 23304
rect 3467 23273 3479 23276
rect 3421 23267 3479 23273
rect 3510 23264 3516 23276
rect 3568 23264 3574 23316
rect 5629 23307 5687 23313
rect 5629 23273 5641 23307
rect 5675 23304 5687 23307
rect 5810 23304 5816 23316
rect 5675 23276 5816 23304
rect 5675 23273 5687 23276
rect 5629 23267 5687 23273
rect 5810 23264 5816 23276
rect 5868 23304 5874 23316
rect 6362 23304 6368 23316
rect 5868 23276 6368 23304
rect 5868 23264 5874 23276
rect 6362 23264 6368 23276
rect 6420 23264 6426 23316
rect 7119 23307 7177 23313
rect 7119 23273 7131 23307
rect 7165 23304 7177 23307
rect 7165 23276 10548 23304
rect 7165 23273 7177 23276
rect 7119 23267 7177 23273
rect 10410 23236 10416 23248
rect 7852 23208 10416 23236
rect 2958 23128 2964 23180
rect 3016 23168 3022 23180
rect 3016 23140 7512 23168
rect 3016 23128 3022 23140
rect 2041 23103 2099 23109
rect 2041 23069 2053 23103
rect 2087 23100 2099 23103
rect 2498 23100 2504 23112
rect 2087 23072 2504 23100
rect 2087 23069 2099 23072
rect 2041 23063 2099 23069
rect 2498 23060 2504 23072
rect 2556 23060 2562 23112
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23100 2743 23103
rect 2774 23100 2780 23112
rect 2731 23072 2780 23100
rect 2731 23069 2743 23072
rect 2685 23063 2743 23069
rect 2774 23060 2780 23072
rect 2832 23060 2838 23112
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23069 7435 23103
rect 7484 23100 7512 23140
rect 7742 23128 7748 23180
rect 7800 23168 7806 23180
rect 7852 23177 7880 23208
rect 10410 23196 10416 23208
rect 10468 23196 10474 23248
rect 10520 23236 10548 23276
rect 10594 23264 10600 23316
rect 10652 23304 10658 23316
rect 10781 23307 10839 23313
rect 10781 23304 10793 23307
rect 10652 23276 10793 23304
rect 10652 23264 10658 23276
rect 10781 23273 10793 23276
rect 10827 23273 10839 23307
rect 10781 23267 10839 23273
rect 10870 23264 10876 23316
rect 10928 23304 10934 23316
rect 16577 23307 16635 23313
rect 10928 23276 11560 23304
rect 10928 23264 10934 23276
rect 11238 23236 11244 23248
rect 10520 23208 11244 23236
rect 11238 23196 11244 23208
rect 11296 23196 11302 23248
rect 7837 23171 7895 23177
rect 7837 23168 7849 23171
rect 7800 23140 7849 23168
rect 7800 23128 7806 23140
rect 7837 23137 7849 23140
rect 7883 23137 7895 23171
rect 7837 23131 7895 23137
rect 7944 23140 9444 23168
rect 7944 23100 7972 23140
rect 8386 23100 8392 23112
rect 7484 23072 7972 23100
rect 8347 23072 8392 23100
rect 7377 23063 7435 23069
rect 4065 23035 4123 23041
rect 4065 23001 4077 23035
rect 4111 23032 4123 23035
rect 4890 23032 4896 23044
rect 4111 23004 4896 23032
rect 4111 23001 4123 23004
rect 4065 22995 4123 23001
rect 4890 22992 4896 23004
rect 4948 23032 4954 23044
rect 5077 23035 5135 23041
rect 5077 23032 5089 23035
rect 4948 23004 5089 23032
rect 4948 22992 4954 23004
rect 5077 23001 5089 23004
rect 5123 23001 5135 23035
rect 6670 23004 7162 23032
rect 5077 22995 5135 23001
rect 2777 22967 2835 22973
rect 2777 22933 2789 22967
rect 2823 22964 2835 22967
rect 3878 22964 3884 22976
rect 2823 22936 3884 22964
rect 2823 22933 2835 22936
rect 2777 22927 2835 22933
rect 3878 22924 3884 22936
rect 3936 22924 3942 22976
rect 4617 22967 4675 22973
rect 4617 22933 4629 22967
rect 4663 22964 4675 22967
rect 5534 22964 5540 22976
rect 4663 22936 5540 22964
rect 4663 22933 4675 22936
rect 4617 22927 4675 22933
rect 5534 22924 5540 22936
rect 5592 22964 5598 22976
rect 6270 22964 6276 22976
rect 5592 22936 6276 22964
rect 5592 22924 5598 22936
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 7134 22964 7162 23004
rect 7190 22992 7196 23044
rect 7248 23032 7254 23044
rect 7392 23032 7420 23063
rect 8386 23060 8392 23072
rect 8444 23060 8450 23112
rect 9416 23109 9444 23140
rect 10594 23128 10600 23180
rect 10652 23168 10658 23180
rect 11425 23171 11483 23177
rect 11425 23168 11437 23171
rect 10652 23140 11437 23168
rect 10652 23128 10658 23140
rect 11425 23137 11437 23140
rect 11471 23137 11483 23171
rect 11532 23168 11560 23276
rect 16577 23273 16589 23307
rect 16623 23304 16635 23307
rect 16666 23304 16672 23316
rect 16623 23276 16672 23304
rect 16623 23273 16635 23276
rect 16577 23267 16635 23273
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 16850 23264 16856 23316
rect 16908 23304 16914 23316
rect 17865 23307 17923 23313
rect 17865 23304 17877 23307
rect 16908 23276 17877 23304
rect 16908 23264 16914 23276
rect 17865 23273 17877 23276
rect 17911 23273 17923 23307
rect 24670 23304 24676 23316
rect 24631 23276 24676 23304
rect 17865 23267 17923 23273
rect 24670 23264 24676 23276
rect 24728 23264 24734 23316
rect 11606 23196 11612 23248
rect 11664 23236 11670 23248
rect 12250 23236 12256 23248
rect 11664 23208 12256 23236
rect 11664 23196 11670 23208
rect 12250 23196 12256 23208
rect 12308 23196 12314 23248
rect 12342 23196 12348 23248
rect 12400 23236 12406 23248
rect 14274 23236 14280 23248
rect 12400 23208 14280 23236
rect 12400 23196 12406 23208
rect 14274 23196 14280 23208
rect 14332 23196 14338 23248
rect 17770 23196 17776 23248
rect 17828 23236 17834 23248
rect 17828 23208 19840 23236
rect 17828 23196 17834 23208
rect 11532 23140 12434 23168
rect 11425 23131 11483 23137
rect 9401 23103 9459 23109
rect 9401 23069 9413 23103
rect 9447 23069 9459 23103
rect 10226 23100 10232 23112
rect 10187 23072 10232 23100
rect 9401 23063 9459 23069
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 10686 23100 10692 23112
rect 10647 23072 10692 23100
rect 10686 23060 10692 23072
rect 10744 23060 10750 23112
rect 12406 23100 12434 23140
rect 13446 23128 13452 23180
rect 13504 23168 13510 23180
rect 13633 23171 13691 23177
rect 13633 23168 13645 23171
rect 13504 23140 13645 23168
rect 13504 23128 13510 23140
rect 13633 23137 13645 23140
rect 13679 23137 13691 23171
rect 13633 23131 13691 23137
rect 15102 23128 15108 23180
rect 15160 23168 15166 23180
rect 15381 23171 15439 23177
rect 15381 23168 15393 23171
rect 15160 23140 15393 23168
rect 15160 23128 15166 23140
rect 15381 23137 15393 23140
rect 15427 23137 15439 23171
rect 15381 23131 15439 23137
rect 16574 23128 16580 23180
rect 16632 23168 16638 23180
rect 17221 23171 17279 23177
rect 17221 23168 17233 23171
rect 16632 23140 17233 23168
rect 16632 23128 16638 23140
rect 17221 23137 17233 23140
rect 17267 23137 17279 23171
rect 19518 23168 19524 23180
rect 19479 23140 19524 23168
rect 17221 23131 17279 23137
rect 19518 23128 19524 23140
rect 19576 23128 19582 23180
rect 19812 23177 19840 23208
rect 19797 23171 19855 23177
rect 19797 23137 19809 23171
rect 19843 23137 19855 23171
rect 19797 23131 19855 23137
rect 14366 23100 14372 23112
rect 12406 23072 13032 23100
rect 14327 23072 14372 23100
rect 7248 23004 7420 23032
rect 8481 23035 8539 23041
rect 7248 22992 7254 23004
rect 8481 23001 8493 23035
rect 8527 23032 8539 23035
rect 8527 23004 10824 23032
rect 8527 23001 8539 23004
rect 8481 22995 8539 23001
rect 8110 22964 8116 22976
rect 7134 22936 8116 22964
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 9490 22964 9496 22976
rect 9451 22936 9496 22964
rect 9490 22924 9496 22936
rect 9548 22924 9554 22976
rect 9582 22924 9588 22976
rect 9640 22964 9646 22976
rect 10137 22967 10195 22973
rect 10137 22964 10149 22967
rect 9640 22936 10149 22964
rect 9640 22924 9646 22936
rect 10137 22933 10149 22936
rect 10183 22933 10195 22967
rect 10796 22964 10824 23004
rect 11238 22992 11244 23044
rect 11296 23032 11302 23044
rect 11422 23032 11428 23044
rect 11296 23004 11428 23032
rect 11296 22992 11302 23004
rect 11422 22992 11428 23004
rect 11480 22992 11486 23044
rect 11514 22992 11520 23044
rect 11572 23032 11578 23044
rect 12069 23035 12127 23041
rect 11572 23004 11617 23032
rect 11572 22992 11578 23004
rect 12069 23001 12081 23035
rect 12115 23032 12127 23035
rect 12158 23032 12164 23044
rect 12115 23004 12164 23032
rect 12115 23001 12127 23004
rect 12069 22995 12127 23001
rect 12158 22992 12164 23004
rect 12216 22992 12222 23044
rect 13004 23041 13032 23072
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 14734 23060 14740 23112
rect 14792 23100 14798 23112
rect 14792 23072 14964 23100
rect 14792 23060 14798 23072
rect 12989 23035 13047 23041
rect 12989 23001 13001 23035
rect 13035 23032 13047 23035
rect 13354 23032 13360 23044
rect 13035 23004 13360 23032
rect 13035 23001 13047 23004
rect 12989 22995 13047 23001
rect 13354 22992 13360 23004
rect 13412 22992 13418 23044
rect 13538 23032 13544 23044
rect 13499 23004 13544 23032
rect 13538 22992 13544 23004
rect 13596 22992 13602 23044
rect 14936 23032 14964 23072
rect 16482 23060 16488 23112
rect 16540 23100 16546 23112
rect 16669 23103 16727 23109
rect 16669 23100 16681 23103
rect 16540 23072 16681 23100
rect 16540 23060 16546 23072
rect 16669 23069 16681 23072
rect 16715 23069 16727 23103
rect 17310 23100 17316 23112
rect 17271 23072 17316 23100
rect 16669 23063 16727 23069
rect 17310 23060 17316 23072
rect 17368 23060 17374 23112
rect 17862 23060 17868 23112
rect 17920 23100 17926 23112
rect 17957 23103 18015 23109
rect 17957 23100 17969 23103
rect 17920 23072 17969 23100
rect 17920 23060 17926 23072
rect 17957 23069 17969 23072
rect 18003 23069 18015 23103
rect 23750 23100 23756 23112
rect 23663 23072 23756 23100
rect 17957 23063 18015 23069
rect 23750 23060 23756 23072
rect 23808 23100 23814 23112
rect 24670 23100 24676 23112
rect 23808 23072 24676 23100
rect 23808 23060 23814 23072
rect 24670 23060 24676 23072
rect 24728 23060 24734 23112
rect 15105 23035 15163 23041
rect 15105 23032 15117 23035
rect 13648 23004 14872 23032
rect 14936 23004 15117 23032
rect 13648 22964 13676 23004
rect 14458 22964 14464 22976
rect 10796 22936 13676 22964
rect 14419 22936 14464 22964
rect 10137 22927 10195 22933
rect 14458 22924 14464 22936
rect 14516 22924 14522 22976
rect 14844 22964 14872 23004
rect 15105 23001 15117 23004
rect 15151 23001 15163 23035
rect 15105 22995 15163 23001
rect 15197 23035 15255 23041
rect 15197 23001 15209 23035
rect 15243 23001 15255 23035
rect 15197 22995 15255 23001
rect 15212 22964 15240 22995
rect 19610 22992 19616 23044
rect 19668 23032 19674 23044
rect 19668 23004 19713 23032
rect 19668 22992 19674 23004
rect 18782 22964 18788 22976
rect 14844 22936 15240 22964
rect 18743 22936 18788 22964
rect 18782 22924 18788 22936
rect 18840 22924 18846 22976
rect 23658 22964 23664 22976
rect 23619 22936 23664 22964
rect 23658 22924 23664 22936
rect 23716 22924 23722 22976
rect 1104 22874 36892 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 36892 22874
rect 1104 22800 36892 22822
rect 1670 22720 1676 22772
rect 1728 22760 1734 22772
rect 1765 22763 1823 22769
rect 1765 22760 1777 22763
rect 1728 22732 1777 22760
rect 1728 22720 1734 22732
rect 1765 22729 1777 22732
rect 1811 22729 1823 22763
rect 1765 22723 1823 22729
rect 3973 22763 4031 22769
rect 3973 22729 3985 22763
rect 4019 22760 4031 22763
rect 4982 22760 4988 22772
rect 4019 22732 4988 22760
rect 4019 22729 4031 22732
rect 3973 22723 4031 22729
rect 4982 22720 4988 22732
rect 5040 22720 5046 22772
rect 7101 22763 7159 22769
rect 7101 22729 7113 22763
rect 7147 22760 7159 22763
rect 8938 22760 8944 22772
rect 7147 22732 8944 22760
rect 7147 22729 7159 22732
rect 7101 22723 7159 22729
rect 8938 22720 8944 22732
rect 8996 22720 9002 22772
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 15933 22763 15991 22769
rect 9548 22732 14964 22760
rect 9548 22720 9554 22732
rect 2774 22692 2780 22704
rect 2240 22664 2780 22692
rect 1578 22624 1584 22636
rect 1539 22596 1584 22624
rect 1578 22584 1584 22596
rect 1636 22584 1642 22636
rect 2240 22633 2268 22664
rect 2774 22652 2780 22664
rect 2832 22652 2838 22704
rect 5994 22692 6000 22704
rect 3726 22664 6000 22692
rect 5994 22652 6000 22664
rect 6052 22652 6058 22704
rect 6270 22652 6276 22704
rect 6328 22692 6334 22704
rect 7282 22692 7288 22704
rect 6328 22664 7288 22692
rect 6328 22652 6334 22664
rect 7282 22652 7288 22664
rect 7340 22652 7346 22704
rect 7929 22695 7987 22701
rect 7929 22661 7941 22695
rect 7975 22692 7987 22695
rect 8018 22692 8024 22704
rect 7975 22664 8024 22692
rect 7975 22661 7987 22664
rect 7929 22655 7987 22661
rect 8018 22652 8024 22664
rect 8076 22652 8082 22704
rect 9858 22692 9864 22704
rect 9154 22664 9864 22692
rect 9858 22652 9864 22664
rect 9916 22652 9922 22704
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 11793 22695 11851 22701
rect 11793 22692 11805 22695
rect 11112 22664 11805 22692
rect 11112 22652 11118 22664
rect 11793 22661 11805 22664
rect 11839 22692 11851 22695
rect 11839 22664 12112 22692
rect 11839 22661 11851 22664
rect 11793 22655 11851 22661
rect 2225 22627 2283 22633
rect 2225 22593 2237 22627
rect 2271 22593 2283 22627
rect 4890 22624 4896 22636
rect 4851 22596 4896 22624
rect 2225 22587 2283 22593
rect 4890 22584 4896 22596
rect 4948 22624 4954 22636
rect 5353 22627 5411 22633
rect 5353 22624 5365 22627
rect 4948 22596 5365 22624
rect 4948 22584 4954 22596
rect 5353 22593 5365 22596
rect 5399 22624 5411 22627
rect 5905 22627 5963 22633
rect 5905 22624 5917 22627
rect 5399 22596 5917 22624
rect 5399 22593 5411 22596
rect 5353 22587 5411 22593
rect 5905 22593 5917 22596
rect 5951 22593 5963 22627
rect 5905 22587 5963 22593
rect 7009 22627 7067 22633
rect 7009 22593 7021 22627
rect 7055 22624 7067 22627
rect 7466 22624 7472 22636
rect 7055 22596 7472 22624
rect 7055 22593 7067 22596
rect 7009 22587 7067 22593
rect 2501 22559 2559 22565
rect 2501 22525 2513 22559
rect 2547 22556 2559 22559
rect 5920 22556 5948 22587
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 10226 22584 10232 22636
rect 10284 22624 10290 22636
rect 10505 22627 10563 22633
rect 10505 22624 10517 22627
rect 10284 22596 10517 22624
rect 10284 22584 10290 22596
rect 10505 22593 10517 22596
rect 10551 22593 10563 22627
rect 10505 22587 10563 22593
rect 7098 22556 7104 22568
rect 2547 22528 5856 22556
rect 5920 22528 7104 22556
rect 2547 22525 2559 22528
rect 2501 22519 2559 22525
rect 4890 22448 4896 22500
rect 4948 22488 4954 22500
rect 5258 22488 5264 22500
rect 4948 22460 5264 22488
rect 4948 22448 4954 22460
rect 5258 22448 5264 22460
rect 5316 22448 5322 22500
rect 5828 22420 5856 22528
rect 7098 22516 7104 22528
rect 7156 22516 7162 22568
rect 7190 22516 7196 22568
rect 7248 22556 7254 22568
rect 7653 22559 7711 22565
rect 7653 22556 7665 22559
rect 7248 22528 7665 22556
rect 7248 22516 7254 22528
rect 7653 22525 7665 22528
rect 7699 22525 7711 22559
rect 10318 22556 10324 22568
rect 7653 22519 7711 22525
rect 7760 22528 10324 22556
rect 6546 22448 6552 22500
rect 6604 22488 6610 22500
rect 7760 22488 7788 22528
rect 10318 22516 10324 22528
rect 10376 22516 10382 22568
rect 10520 22556 10548 22587
rect 10594 22584 10600 22636
rect 10652 22624 10658 22636
rect 11885 22627 11943 22633
rect 10652 22614 11100 22624
rect 11149 22617 11207 22623
rect 11149 22614 11161 22617
rect 10652 22596 11161 22614
rect 10652 22584 10658 22596
rect 11072 22586 11161 22596
rect 11149 22583 11161 22586
rect 11195 22583 11207 22617
rect 11885 22593 11897 22627
rect 11931 22624 11943 22627
rect 11974 22624 11980 22636
rect 11931 22596 11980 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 11974 22584 11980 22596
rect 12032 22584 12038 22636
rect 11149 22577 11207 22583
rect 10870 22556 10876 22568
rect 10520 22528 10876 22556
rect 10870 22516 10876 22528
rect 10928 22516 10934 22568
rect 12084 22556 12112 22664
rect 12250 22652 12256 22704
rect 12308 22692 12314 22704
rect 12529 22695 12587 22701
rect 12529 22692 12541 22695
rect 12308 22664 12541 22692
rect 12308 22652 12314 22664
rect 12529 22661 12541 22664
rect 12575 22661 12587 22695
rect 12529 22655 12587 22661
rect 13354 22652 13360 22704
rect 13412 22692 13418 22704
rect 14277 22695 14335 22701
rect 14277 22692 14289 22695
rect 13412 22664 14289 22692
rect 13412 22652 13418 22664
rect 14277 22661 14289 22664
rect 14323 22661 14335 22695
rect 14277 22655 14335 22661
rect 14458 22652 14464 22704
rect 14516 22692 14522 22704
rect 14829 22695 14887 22701
rect 14829 22692 14841 22695
rect 14516 22664 14841 22692
rect 14516 22652 14522 22664
rect 14829 22661 14841 22664
rect 14875 22661 14887 22695
rect 14936 22692 14964 22732
rect 15933 22729 15945 22763
rect 15979 22760 15991 22763
rect 16206 22760 16212 22772
rect 15979 22732 16212 22760
rect 15979 22729 15991 22732
rect 15933 22723 15991 22729
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 18046 22720 18052 22772
rect 18104 22760 18110 22772
rect 18141 22763 18199 22769
rect 18141 22760 18153 22763
rect 18104 22732 18153 22760
rect 18104 22720 18110 22732
rect 18141 22729 18153 22732
rect 18187 22729 18199 22763
rect 18141 22723 18199 22729
rect 17037 22695 17095 22701
rect 17037 22692 17049 22695
rect 14936 22664 17049 22692
rect 14829 22655 14887 22661
rect 17037 22661 17049 22664
rect 17083 22661 17095 22695
rect 17037 22655 17095 22661
rect 17589 22695 17647 22701
rect 17589 22661 17601 22695
rect 17635 22692 17647 22695
rect 21174 22692 21180 22704
rect 17635 22664 21180 22692
rect 17635 22661 17647 22664
rect 17589 22655 17647 22661
rect 13722 22624 13728 22636
rect 13683 22596 13728 22624
rect 13722 22584 13728 22596
rect 13780 22584 13786 22636
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 12084 22528 12449 22556
rect 12437 22525 12449 22528
rect 12483 22525 12495 22559
rect 14918 22556 14924 22568
rect 14879 22528 14924 22556
rect 12437 22519 12495 22525
rect 14918 22516 14924 22528
rect 14976 22516 14982 22568
rect 16945 22559 17003 22565
rect 16945 22525 16957 22559
rect 16991 22556 17003 22559
rect 17954 22556 17960 22568
rect 16991 22528 17960 22556
rect 16991 22525 17003 22528
rect 16945 22519 17003 22525
rect 17954 22516 17960 22528
rect 18012 22516 18018 22568
rect 6604 22460 7788 22488
rect 8956 22460 9674 22488
rect 6604 22448 6610 22460
rect 7374 22420 7380 22432
rect 5828 22392 7380 22420
rect 7374 22380 7380 22392
rect 7432 22420 7438 22432
rect 7926 22420 7932 22432
rect 7432 22392 7932 22420
rect 7432 22380 7438 22392
rect 7926 22380 7932 22392
rect 7984 22380 7990 22432
rect 8294 22380 8300 22432
rect 8352 22420 8358 22432
rect 8956 22420 8984 22460
rect 8352 22392 8984 22420
rect 8352 22380 8358 22392
rect 9030 22380 9036 22432
rect 9088 22420 9094 22432
rect 9401 22423 9459 22429
rect 9401 22420 9413 22423
rect 9088 22392 9413 22420
rect 9088 22380 9094 22392
rect 9401 22389 9413 22392
rect 9447 22389 9459 22423
rect 9646 22420 9674 22460
rect 9766 22448 9772 22500
rect 9824 22488 9830 22500
rect 10594 22488 10600 22500
rect 9824 22460 10600 22488
rect 9824 22448 9830 22460
rect 10594 22448 10600 22460
rect 10652 22448 10658 22500
rect 12989 22491 13047 22497
rect 12989 22457 13001 22491
rect 13035 22488 13047 22491
rect 13170 22488 13176 22500
rect 13035 22460 13176 22488
rect 13035 22457 13047 22460
rect 12989 22451 13047 22457
rect 13170 22448 13176 22460
rect 13228 22448 13234 22500
rect 13354 22448 13360 22500
rect 13412 22488 13418 22500
rect 13722 22488 13728 22500
rect 13412 22460 13728 22488
rect 13412 22448 13418 22460
rect 13722 22448 13728 22460
rect 13780 22448 13786 22500
rect 15102 22448 15108 22500
rect 15160 22488 15166 22500
rect 18064 22488 18092 22664
rect 21174 22652 21180 22664
rect 21232 22652 21238 22704
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22624 18291 22627
rect 18693 22627 18751 22633
rect 18693 22624 18705 22627
rect 18279 22596 18705 22624
rect 18279 22593 18291 22596
rect 18233 22587 18291 22593
rect 18693 22593 18705 22596
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22624 19763 22627
rect 20254 22624 20260 22636
rect 19751 22596 20260 22624
rect 19751 22593 19763 22596
rect 19705 22587 19763 22593
rect 15160 22460 18092 22488
rect 15160 22448 15166 22460
rect 10413 22423 10471 22429
rect 10413 22420 10425 22423
rect 9646 22392 10425 22420
rect 9401 22383 9459 22389
rect 10413 22389 10425 22392
rect 10459 22389 10471 22423
rect 11054 22420 11060 22432
rect 11015 22392 11060 22420
rect 10413 22383 10471 22389
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 11146 22380 11152 22432
rect 11204 22420 11210 22432
rect 12342 22420 12348 22432
rect 11204 22392 12348 22420
rect 11204 22380 11210 22392
rect 12342 22380 12348 22392
rect 12400 22380 12406 22432
rect 13078 22380 13084 22432
rect 13136 22420 13142 22432
rect 13633 22423 13691 22429
rect 13633 22420 13645 22423
rect 13136 22392 13645 22420
rect 13136 22380 13142 22392
rect 13633 22389 13645 22392
rect 13679 22389 13691 22423
rect 13633 22383 13691 22389
rect 14918 22380 14924 22432
rect 14976 22420 14982 22432
rect 15470 22420 15476 22432
rect 14976 22392 15476 22420
rect 14976 22380 14982 22392
rect 15470 22380 15476 22392
rect 15528 22380 15534 22432
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 18248 22420 18276 22587
rect 20254 22584 20260 22596
rect 20312 22584 20318 22636
rect 24854 22584 24860 22636
rect 24912 22624 24918 22636
rect 28629 22627 28687 22633
rect 28629 22624 28641 22627
rect 24912 22596 28641 22624
rect 24912 22584 24918 22596
rect 28629 22593 28641 22596
rect 28675 22593 28687 22627
rect 28629 22587 28687 22593
rect 28721 22627 28779 22633
rect 28721 22593 28733 22627
rect 28767 22624 28779 22627
rect 36081 22627 36139 22633
rect 36081 22624 36093 22627
rect 28767 22596 36093 22624
rect 28767 22593 28779 22596
rect 28721 22587 28779 22593
rect 36081 22593 36093 22596
rect 36127 22593 36139 22627
rect 36081 22587 36139 22593
rect 28644 22556 28672 22587
rect 29273 22559 29331 22565
rect 29273 22556 29285 22559
rect 28644 22528 29285 22556
rect 29273 22525 29285 22528
rect 29319 22525 29331 22559
rect 29273 22519 29331 22525
rect 36262 22488 36268 22500
rect 36223 22460 36268 22488
rect 36262 22448 36268 22460
rect 36320 22448 36326 22500
rect 19610 22420 19616 22432
rect 16816 22392 18276 22420
rect 19571 22392 19616 22420
rect 16816 22380 16822 22392
rect 19610 22380 19616 22392
rect 19668 22380 19674 22432
rect 20254 22420 20260 22432
rect 20215 22392 20260 22420
rect 20254 22380 20260 22392
rect 20312 22380 20318 22432
rect 1104 22330 36892 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 36892 22330
rect 1104 22256 36892 22278
rect 4236 22219 4294 22225
rect 4236 22185 4248 22219
rect 4282 22216 4294 22219
rect 4982 22216 4988 22228
rect 4282 22188 4988 22216
rect 4282 22185 4294 22188
rect 4236 22179 4294 22185
rect 4982 22176 4988 22188
rect 5040 22176 5046 22228
rect 7098 22176 7104 22228
rect 7156 22216 7162 22228
rect 7156 22188 7880 22216
rect 7156 22176 7162 22188
rect 5276 22120 6224 22148
rect 3234 22040 3240 22092
rect 3292 22080 3298 22092
rect 5276 22080 5304 22120
rect 3292 22052 5304 22080
rect 3292 22040 3298 22052
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 2314 22012 2320 22024
rect 1903 21984 2320 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 2314 21972 2320 21984
rect 2372 21972 2378 22024
rect 2774 21972 2780 22024
rect 2832 22012 2838 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 2832 21984 3985 22012
rect 2832 21972 2838 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 5258 21904 5264 21956
rect 5316 21904 5322 21956
rect 6196 21944 6224 22120
rect 6273 22083 6331 22089
rect 6273 22049 6285 22083
rect 6319 22080 6331 22083
rect 7190 22080 7196 22092
rect 6319 22052 7196 22080
rect 6319 22049 6331 22052
rect 6273 22043 6331 22049
rect 7190 22040 7196 22052
rect 7248 22040 7254 22092
rect 7852 22080 7880 22188
rect 7926 22176 7932 22228
rect 7984 22216 7990 22228
rect 8021 22219 8079 22225
rect 8021 22216 8033 22219
rect 7984 22188 8033 22216
rect 7984 22176 7990 22188
rect 8021 22185 8033 22188
rect 8067 22185 8079 22219
rect 8021 22179 8079 22185
rect 9490 22176 9496 22228
rect 9548 22216 9554 22228
rect 11146 22216 11152 22228
rect 9548 22188 11152 22216
rect 9548 22176 9554 22188
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 11241 22219 11299 22225
rect 11241 22185 11253 22219
rect 11287 22216 11299 22219
rect 11514 22216 11520 22228
rect 11287 22188 11520 22216
rect 11287 22185 11299 22188
rect 11241 22179 11299 22185
rect 11514 22176 11520 22188
rect 11572 22176 11578 22228
rect 12529 22219 12587 22225
rect 12529 22185 12541 22219
rect 12575 22216 12587 22219
rect 13538 22216 13544 22228
rect 12575 22188 13544 22216
rect 12575 22185 12587 22188
rect 12529 22179 12587 22185
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 14918 22216 14924 22228
rect 13832 22188 14924 22216
rect 9122 22108 9128 22160
rect 9180 22148 9186 22160
rect 9674 22148 9680 22160
rect 9180 22120 9680 22148
rect 9180 22108 9186 22120
rect 9674 22108 9680 22120
rect 9732 22108 9738 22160
rect 9766 22108 9772 22160
rect 9824 22108 9830 22160
rect 9876 22120 11836 22148
rect 9784 22080 9812 22108
rect 7852 22052 9812 22080
rect 7650 21972 7656 22024
rect 7708 21972 7714 22024
rect 8110 21972 8116 22024
rect 8168 22012 8174 22024
rect 9214 22012 9220 22024
rect 8168 21984 9220 22012
rect 8168 21972 8174 21984
rect 9214 21972 9220 21984
rect 9272 21972 9278 22024
rect 9416 22021 9444 22052
rect 9401 22015 9459 22021
rect 9401 21981 9413 22015
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 9876 22022 9904 22120
rect 10060 22080 10272 22092
rect 10597 22083 10655 22089
rect 10060 22064 10364 22080
rect 10060 22031 10088 22064
rect 10244 22052 10364 22064
rect 9692 22012 9904 22022
rect 9548 21994 9904 22012
rect 10045 22025 10103 22031
rect 9548 21984 9720 21994
rect 10045 21991 10057 22025
rect 10091 21991 10103 22025
rect 10045 21985 10103 21991
rect 9548 21972 9554 21984
rect 6546 21944 6552 21956
rect 6196 21916 6552 21944
rect 6546 21904 6552 21916
rect 6604 21904 6610 21956
rect 9416 21916 9674 21944
rect 9416 21888 9444 21916
rect 1670 21876 1676 21888
rect 1631 21848 1676 21876
rect 1670 21836 1676 21848
rect 1728 21836 1734 21888
rect 2869 21879 2927 21885
rect 2869 21845 2881 21879
rect 2915 21876 2927 21879
rect 3050 21876 3056 21888
rect 2915 21848 3056 21876
rect 2915 21845 2927 21848
rect 2869 21839 2927 21845
rect 3050 21836 3056 21848
rect 3108 21836 3114 21888
rect 3234 21836 3240 21888
rect 3292 21876 3298 21888
rect 3329 21879 3387 21885
rect 3329 21876 3341 21879
rect 3292 21848 3341 21876
rect 3292 21836 3298 21848
rect 3329 21845 3341 21848
rect 3375 21845 3387 21879
rect 3329 21839 3387 21845
rect 4982 21836 4988 21888
rect 5040 21876 5046 21888
rect 5721 21879 5779 21885
rect 5721 21876 5733 21879
rect 5040 21848 5733 21876
rect 5040 21836 5046 21848
rect 5721 21845 5733 21848
rect 5767 21845 5779 21879
rect 5721 21839 5779 21845
rect 6454 21836 6460 21888
rect 6512 21876 6518 21888
rect 8570 21876 8576 21888
rect 6512 21848 8576 21876
rect 6512 21836 6518 21848
rect 8570 21836 8576 21848
rect 8628 21836 8634 21888
rect 9306 21876 9312 21888
rect 9267 21848 9312 21876
rect 9306 21836 9312 21848
rect 9364 21836 9370 21888
rect 9398 21836 9404 21888
rect 9456 21836 9462 21888
rect 9646 21876 9674 21916
rect 9766 21904 9772 21956
rect 9824 21904 9830 21956
rect 10336 21944 10364 22052
rect 10597 22049 10609 22083
rect 10643 22080 10655 22083
rect 10778 22080 10784 22092
rect 10643 22052 10784 22080
rect 10643 22049 10655 22052
rect 10597 22043 10655 22049
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 10410 21972 10416 22024
rect 10468 22006 10474 22024
rect 10505 22015 10563 22021
rect 10505 22006 10517 22015
rect 10468 21981 10517 22006
rect 10551 21981 10563 22015
rect 10468 21978 10563 21981
rect 10468 21972 10474 21978
rect 10505 21975 10563 21978
rect 11149 22015 11207 22021
rect 11149 21981 11161 22015
rect 11195 22012 11207 22015
rect 11238 22012 11244 22024
rect 11195 21984 11244 22012
rect 11195 21981 11207 21984
rect 11149 21975 11207 21981
rect 11238 21972 11244 21984
rect 11296 21972 11302 22024
rect 11808 22021 11836 22120
rect 13541 22083 13599 22089
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 13630 22080 13636 22092
rect 13587 22052 13636 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 13630 22040 13636 22052
rect 13688 22040 13694 22092
rect 13722 22040 13728 22092
rect 13780 22080 13786 22092
rect 13832 22080 13860 22188
rect 14918 22176 14924 22188
rect 14976 22176 14982 22228
rect 15470 22176 15476 22228
rect 15528 22216 15534 22228
rect 19610 22216 19616 22228
rect 15528 22188 19616 22216
rect 15528 22176 15534 22188
rect 19610 22176 19616 22188
rect 19668 22176 19674 22228
rect 18046 22148 18052 22160
rect 13780 22052 13860 22080
rect 14292 22120 18052 22148
rect 13780 22040 13786 22052
rect 12437 22025 12495 22031
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 21981 11851 22015
rect 11793 21975 11851 21981
rect 10870 21944 10876 21956
rect 10336 21916 10876 21944
rect 10870 21904 10876 21916
rect 10928 21904 10934 21956
rect 11808 21944 11836 21975
rect 11974 21972 11980 22024
rect 12032 22012 12038 22024
rect 12437 22022 12449 22025
rect 12268 22012 12449 22022
rect 12032 21994 12449 22012
rect 12032 21984 12296 21994
rect 12437 21991 12449 21994
rect 12483 21991 12495 22025
rect 12437 21985 12495 21991
rect 13081 22015 13139 22021
rect 12032 21972 12038 21984
rect 13081 21981 13093 22015
rect 13127 22012 13139 22015
rect 14090 22012 14096 22024
rect 13127 21984 14096 22012
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 14292 21944 14320 22120
rect 18046 22108 18052 22120
rect 18104 22148 18110 22160
rect 18598 22148 18604 22160
rect 18104 22120 18604 22148
rect 18104 22108 18110 22120
rect 18598 22108 18604 22120
rect 18656 22108 18662 22160
rect 14458 22080 14464 22092
rect 14419 22052 14464 22080
rect 14458 22040 14464 22052
rect 14516 22040 14522 22092
rect 14918 22080 14924 22092
rect 14879 22052 14924 22080
rect 14918 22040 14924 22052
rect 14976 22040 14982 22092
rect 15194 22040 15200 22092
rect 15252 22080 15258 22092
rect 15252 22052 15516 22080
rect 15252 22040 15258 22052
rect 15488 22021 15516 22052
rect 15930 22040 15936 22092
rect 15988 22080 15994 22092
rect 16500 22089 16620 22092
rect 16500 22083 16635 22089
rect 16500 22080 16589 22083
rect 15988 22064 16589 22080
rect 15988 22052 16528 22064
rect 15988 22040 15994 22052
rect 16577 22049 16589 22064
rect 16623 22049 16635 22083
rect 16577 22043 16635 22049
rect 15473 22015 15531 22021
rect 15473 21981 15485 22015
rect 15519 22012 15531 22015
rect 16206 22012 16212 22024
rect 15519 21984 16212 22012
rect 15519 21981 15531 21984
rect 15473 21975 15531 21981
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 19981 22015 20039 22021
rect 19981 21981 19993 22015
rect 20027 22012 20039 22015
rect 20714 22012 20720 22024
rect 20027 21984 20720 22012
rect 20027 21981 20039 21984
rect 19981 21975 20039 21981
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 26329 22015 26387 22021
rect 26329 21981 26341 22015
rect 26375 22012 26387 22015
rect 35894 22012 35900 22024
rect 26375 21984 35900 22012
rect 26375 21981 26387 21984
rect 26329 21975 26387 21981
rect 35894 21972 35900 21984
rect 35952 21972 35958 22024
rect 11808 21916 14320 21944
rect 14829 21947 14887 21953
rect 14829 21913 14841 21947
rect 14875 21944 14887 21947
rect 15194 21944 15200 21956
rect 14875 21916 15200 21944
rect 14875 21913 14887 21916
rect 14829 21907 14887 21913
rect 15194 21904 15200 21916
rect 15252 21904 15258 21956
rect 17126 21944 17132 21956
rect 17087 21916 17132 21944
rect 17126 21904 17132 21916
rect 17184 21904 17190 21956
rect 17218 21904 17224 21956
rect 17276 21944 17282 21956
rect 18141 21947 18199 21953
rect 18141 21944 18153 21947
rect 17276 21916 18153 21944
rect 17276 21904 17282 21916
rect 18141 21913 18153 21916
rect 18187 21913 18199 21947
rect 18141 21907 18199 21913
rect 18230 21904 18236 21956
rect 18288 21944 18294 21956
rect 18785 21947 18843 21953
rect 18288 21916 18333 21944
rect 18288 21904 18294 21916
rect 18785 21913 18797 21947
rect 18831 21944 18843 21947
rect 19242 21944 19248 21956
rect 18831 21916 19248 21944
rect 18831 21913 18843 21916
rect 18785 21907 18843 21913
rect 9784 21876 9812 21904
rect 9646 21848 9812 21876
rect 9953 21879 10011 21885
rect 9953 21845 9965 21879
rect 9999 21876 10011 21879
rect 10042 21876 10048 21888
rect 9999 21848 10048 21876
rect 9999 21845 10011 21848
rect 9953 21839 10011 21845
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 11885 21879 11943 21885
rect 11885 21845 11897 21879
rect 11931 21876 11943 21879
rect 12894 21876 12900 21888
rect 11931 21848 12900 21876
rect 11931 21845 11943 21848
rect 11885 21839 11943 21845
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 15562 21876 15568 21888
rect 15523 21848 15568 21876
rect 15562 21836 15568 21848
rect 15620 21836 15626 21888
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 18800 21876 18828 21907
rect 19242 21904 19248 21916
rect 19300 21904 19306 21956
rect 22002 21944 22008 21956
rect 20180 21916 22008 21944
rect 20180 21885 20208 21916
rect 22002 21904 22008 21916
rect 22060 21904 22066 21956
rect 18012 21848 18828 21876
rect 20165 21879 20223 21885
rect 18012 21836 18018 21848
rect 20165 21845 20177 21879
rect 20211 21845 20223 21879
rect 20714 21876 20720 21888
rect 20675 21848 20720 21876
rect 20165 21839 20223 21845
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 21818 21876 21824 21888
rect 21324 21848 21824 21876
rect 21324 21836 21330 21848
rect 21818 21836 21824 21848
rect 21876 21876 21882 21888
rect 26237 21879 26295 21885
rect 26237 21876 26249 21879
rect 21876 21848 26249 21876
rect 21876 21836 21882 21848
rect 26237 21845 26249 21848
rect 26283 21845 26295 21879
rect 26237 21839 26295 21845
rect 1104 21786 36892 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 36892 21786
rect 1104 21712 36892 21734
rect 6822 21672 6828 21684
rect 6783 21644 6828 21672
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 10045 21675 10103 21681
rect 10045 21672 10057 21675
rect 7392 21644 10057 21672
rect 7392 21604 7420 21644
rect 10045 21641 10057 21644
rect 10091 21641 10103 21675
rect 10045 21635 10103 21641
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 11977 21675 12035 21681
rect 11977 21672 11989 21675
rect 11940 21644 11989 21672
rect 11940 21632 11946 21644
rect 11977 21641 11989 21644
rect 12023 21641 12035 21675
rect 12618 21672 12624 21684
rect 12579 21644 12624 21672
rect 11977 21635 12035 21641
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 16945 21675 17003 21681
rect 12728 21644 14596 21672
rect 7558 21604 7564 21616
rect 4830 21576 7420 21604
rect 7519 21576 7564 21604
rect 7558 21564 7564 21576
rect 7616 21564 7622 21616
rect 10410 21604 10416 21616
rect 8786 21576 10416 21604
rect 10410 21564 10416 21576
rect 10468 21564 10474 21616
rect 10686 21564 10692 21616
rect 10744 21604 10750 21616
rect 10744 21576 11008 21604
rect 10744 21564 10750 21576
rect 1854 21536 1860 21548
rect 1815 21508 1860 21536
rect 1854 21496 1860 21508
rect 1912 21496 1918 21548
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 10137 21539 10195 21545
rect 8996 21508 9444 21536
rect 8996 21496 9002 21508
rect 9416 21480 9444 21508
rect 10137 21505 10149 21539
rect 10183 21536 10195 21539
rect 10594 21536 10600 21548
rect 10183 21508 10600 21536
rect 10183 21505 10195 21508
rect 10137 21499 10195 21505
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21536 10839 21539
rect 10870 21536 10876 21548
rect 10827 21508 10876 21536
rect 10827 21505 10839 21508
rect 10781 21499 10839 21505
rect 10870 21496 10876 21508
rect 10928 21496 10934 21548
rect 10980 21536 11008 21576
rect 11146 21564 11152 21616
rect 11204 21604 11210 21616
rect 12728 21604 12756 21644
rect 11204 21576 12756 21604
rect 11204 21564 11210 21576
rect 13630 21564 13636 21616
rect 13688 21604 13694 21616
rect 13725 21607 13783 21613
rect 13725 21604 13737 21607
rect 13688 21576 13737 21604
rect 13688 21564 13694 21576
rect 13725 21573 13737 21576
rect 13771 21573 13783 21607
rect 13725 21567 13783 21573
rect 14182 21564 14188 21616
rect 14240 21604 14246 21616
rect 14458 21604 14464 21616
rect 14240 21576 14464 21604
rect 14240 21564 14246 21576
rect 14458 21564 14464 21576
rect 14516 21564 14522 21616
rect 14568 21613 14596 21644
rect 16945 21641 16957 21675
rect 16991 21672 17003 21675
rect 17034 21672 17040 21684
rect 16991 21644 17040 21672
rect 16991 21641 17003 21644
rect 16945 21635 17003 21641
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 14553 21607 14611 21613
rect 14553 21573 14565 21607
rect 14599 21573 14611 21607
rect 15102 21604 15108 21616
rect 15063 21576 15108 21604
rect 14553 21567 14611 21573
rect 15102 21564 15108 21576
rect 15160 21564 15166 21616
rect 15378 21564 15384 21616
rect 15436 21604 15442 21616
rect 15565 21607 15623 21613
rect 15565 21604 15577 21607
rect 15436 21576 15577 21604
rect 15436 21564 15442 21576
rect 15565 21573 15577 21576
rect 15611 21573 15623 21607
rect 16114 21604 16120 21616
rect 16075 21576 16120 21604
rect 15565 21567 15623 21573
rect 16114 21564 16120 21576
rect 16172 21564 16178 21616
rect 16206 21564 16212 21616
rect 16264 21604 16270 21616
rect 18141 21607 18199 21613
rect 18141 21604 18153 21607
rect 16264 21576 18153 21604
rect 16264 21564 16270 21576
rect 18141 21573 18153 21576
rect 18187 21573 18199 21607
rect 18141 21567 18199 21573
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 10980 21508 12081 21536
rect 12069 21505 12081 21508
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 12526 21496 12532 21548
rect 12584 21536 12590 21548
rect 12713 21539 12771 21545
rect 12713 21536 12725 21539
rect 12584 21508 12725 21536
rect 12584 21496 12590 21508
rect 12713 21505 12725 21508
rect 12759 21505 12771 21539
rect 16850 21536 16856 21548
rect 16811 21508 16856 21536
rect 12713 21499 12771 21505
rect 16850 21496 16856 21508
rect 16908 21496 16914 21548
rect 35621 21539 35679 21545
rect 35621 21505 35633 21539
rect 35667 21536 35679 21539
rect 36262 21536 36268 21548
rect 35667 21508 36268 21536
rect 35667 21505 35679 21508
rect 35621 21499 35679 21505
rect 36262 21496 36268 21508
rect 36320 21496 36326 21548
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 3329 21471 3387 21477
rect 3329 21468 3341 21471
rect 2832 21440 3341 21468
rect 2832 21428 2838 21440
rect 3329 21437 3341 21440
rect 3375 21437 3387 21471
rect 3602 21468 3608 21480
rect 3563 21440 3608 21468
rect 3329 21431 3387 21437
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21468 5411 21471
rect 5442 21468 5448 21480
rect 5399 21440 5448 21468
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 5442 21428 5448 21440
rect 5500 21428 5506 21480
rect 5997 21471 6055 21477
rect 5997 21437 6009 21471
rect 6043 21468 6055 21471
rect 6822 21468 6828 21480
rect 6043 21440 6828 21468
rect 6043 21437 6055 21440
rect 5997 21431 6055 21437
rect 6822 21428 6828 21440
rect 6880 21428 6886 21480
rect 7190 21428 7196 21480
rect 7248 21468 7254 21480
rect 7285 21471 7343 21477
rect 7285 21468 7297 21471
rect 7248 21440 7297 21468
rect 7248 21428 7254 21440
rect 7285 21437 7297 21440
rect 7331 21437 7343 21471
rect 7285 21431 7343 21437
rect 8754 21428 8760 21480
rect 8812 21468 8818 21480
rect 9030 21468 9036 21480
rect 8812 21440 9036 21468
rect 8812 21428 8818 21440
rect 9030 21428 9036 21440
rect 9088 21468 9094 21480
rect 9309 21471 9367 21477
rect 9309 21468 9321 21471
rect 9088 21440 9321 21468
rect 9088 21428 9094 21440
rect 9309 21437 9321 21440
rect 9355 21437 9367 21471
rect 9309 21431 9367 21437
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 13541 21471 13599 21477
rect 9456 21440 12388 21468
rect 9456 21428 9462 21440
rect 12360 21412 12388 21440
rect 13541 21437 13553 21471
rect 13587 21437 13599 21471
rect 13541 21431 13599 21437
rect 4614 21360 4620 21412
rect 4672 21400 4678 21412
rect 4672 21372 6868 21400
rect 4672 21360 4678 21372
rect 1670 21332 1676 21344
rect 1631 21304 1676 21332
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 2866 21332 2872 21344
rect 2827 21304 2872 21332
rect 2866 21292 2872 21304
rect 2924 21292 2930 21344
rect 6840 21332 6868 21372
rect 8662 21360 8668 21412
rect 8720 21400 8726 21412
rect 8720 21372 10824 21400
rect 8720 21360 8726 21372
rect 10689 21335 10747 21341
rect 10689 21332 10701 21335
rect 6840 21304 10701 21332
rect 10689 21301 10701 21304
rect 10735 21301 10747 21335
rect 10796 21332 10824 21372
rect 12342 21360 12348 21412
rect 12400 21400 12406 21412
rect 13556 21400 13584 21431
rect 13722 21428 13728 21480
rect 13780 21468 13786 21480
rect 13817 21471 13875 21477
rect 13817 21468 13829 21471
rect 13780 21440 13829 21468
rect 13780 21428 13786 21440
rect 13817 21437 13829 21440
rect 13863 21437 13875 21471
rect 13817 21431 13875 21437
rect 14274 21428 14280 21480
rect 14332 21468 14338 21480
rect 14458 21468 14464 21480
rect 14332 21440 14464 21468
rect 14332 21428 14338 21440
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 16209 21471 16267 21477
rect 16209 21437 16221 21471
rect 16255 21468 16267 21471
rect 19426 21468 19432 21480
rect 16255 21440 19432 21468
rect 16255 21437 16267 21440
rect 16209 21431 16267 21437
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 13998 21400 14004 21412
rect 12400 21372 13492 21400
rect 13556 21372 14004 21400
rect 12400 21360 12406 21372
rect 12710 21332 12716 21344
rect 10796 21304 12716 21332
rect 10689 21295 10747 21301
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 13464 21332 13492 21372
rect 13998 21360 14004 21372
rect 14056 21400 14062 21412
rect 14642 21400 14648 21412
rect 14056 21372 14648 21400
rect 14056 21360 14062 21372
rect 14642 21360 14648 21372
rect 14700 21360 14706 21412
rect 15010 21360 15016 21412
rect 15068 21400 15074 21412
rect 18693 21403 18751 21409
rect 18693 21400 18705 21403
rect 15068 21372 18705 21400
rect 15068 21360 15074 21372
rect 18693 21369 18705 21372
rect 18739 21369 18751 21403
rect 18693 21363 18751 21369
rect 18782 21360 18788 21412
rect 18840 21400 18846 21412
rect 21910 21400 21916 21412
rect 18840 21372 21916 21400
rect 18840 21360 18846 21372
rect 21910 21360 21916 21372
rect 21968 21400 21974 21412
rect 35986 21400 35992 21412
rect 21968 21372 35992 21400
rect 21968 21360 21974 21372
rect 35986 21360 35992 21372
rect 36044 21360 36050 21412
rect 16850 21332 16856 21344
rect 13464 21304 16856 21332
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 17586 21332 17592 21344
rect 17547 21304 17592 21332
rect 17586 21292 17592 21304
rect 17644 21332 17650 21344
rect 17862 21332 17868 21344
rect 17644 21304 17868 21332
rect 17644 21292 17650 21304
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 36170 21332 36176 21344
rect 36131 21304 36176 21332
rect 36170 21292 36176 21304
rect 36228 21292 36234 21344
rect 1104 21242 36892 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 36892 21242
rect 1104 21168 36892 21190
rect 2133 21131 2191 21137
rect 2133 21097 2145 21131
rect 2179 21128 2191 21131
rect 2774 21128 2780 21140
rect 2179 21100 2780 21128
rect 2179 21097 2191 21100
rect 2133 21091 2191 21097
rect 2774 21088 2780 21100
rect 2832 21088 2838 21140
rect 2866 21088 2872 21140
rect 2924 21128 2930 21140
rect 8386 21128 8392 21140
rect 2924 21100 8392 21128
rect 2924 21088 2930 21100
rect 8386 21088 8392 21100
rect 8444 21128 8450 21140
rect 9122 21128 9128 21140
rect 8444 21100 9128 21128
rect 8444 21088 8450 21100
rect 9122 21088 9128 21100
rect 9180 21088 9186 21140
rect 10962 21128 10968 21140
rect 10923 21100 10968 21128
rect 10962 21088 10968 21100
rect 11020 21088 11026 21140
rect 12250 21128 12256 21140
rect 12211 21100 12256 21128
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 15010 21128 15016 21140
rect 12360 21100 15016 21128
rect 8754 21020 8760 21072
rect 8812 21060 8818 21072
rect 9398 21060 9404 21072
rect 8812 21032 9404 21060
rect 8812 21020 8818 21032
rect 9398 21020 9404 21032
rect 9456 21020 9462 21072
rect 9677 21063 9735 21069
rect 9677 21029 9689 21063
rect 9723 21060 9735 21063
rect 11146 21060 11152 21072
rect 9723 21032 11152 21060
rect 9723 21029 9735 21032
rect 9677 21023 9735 21029
rect 11146 21020 11152 21032
rect 11204 21020 11210 21072
rect 4341 20995 4399 21001
rect 4341 20961 4353 20995
rect 4387 20992 4399 20995
rect 4982 20992 4988 21004
rect 4387 20964 4988 20992
rect 4387 20961 4399 20964
rect 4341 20955 4399 20961
rect 4982 20952 4988 20964
rect 5040 20952 5046 21004
rect 5074 20952 5080 21004
rect 5132 20992 5138 21004
rect 6089 20995 6147 21001
rect 6089 20992 6101 20995
rect 5132 20964 6101 20992
rect 5132 20952 5138 20964
rect 6089 20961 6101 20964
rect 6135 20992 6147 20995
rect 6454 20992 6460 21004
rect 6135 20964 6460 20992
rect 6135 20961 6147 20964
rect 6089 20955 6147 20961
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 6822 20952 6828 21004
rect 6880 20992 6886 21004
rect 8938 20992 8944 21004
rect 6880 20964 8944 20992
rect 6880 20952 6886 20964
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 9490 20952 9496 21004
rect 9548 20992 9554 21004
rect 10321 20995 10379 21001
rect 10321 20992 10333 20995
rect 9548 20964 10333 20992
rect 9548 20952 9554 20964
rect 10321 20961 10333 20964
rect 10367 20961 10379 20995
rect 12360 20992 12388 21100
rect 15010 21088 15016 21100
rect 15068 21088 15074 21140
rect 16945 21131 17003 21137
rect 16945 21097 16957 21131
rect 16991 21128 17003 21131
rect 18230 21128 18236 21140
rect 16991 21100 18236 21128
rect 16991 21097 17003 21100
rect 16945 21091 17003 21097
rect 18230 21088 18236 21100
rect 18288 21088 18294 21140
rect 18693 21131 18751 21137
rect 18693 21097 18705 21131
rect 18739 21128 18751 21131
rect 18782 21128 18788 21140
rect 18739 21100 18788 21128
rect 18739 21097 18751 21100
rect 18693 21091 18751 21097
rect 18782 21088 18788 21100
rect 18840 21088 18846 21140
rect 13449 21063 13507 21069
rect 13449 21029 13461 21063
rect 13495 21060 13507 21063
rect 13495 21032 15332 21060
rect 13495 21029 13507 21032
rect 13449 21023 13507 21029
rect 10321 20955 10379 20961
rect 10888 20964 12388 20992
rect 2774 20884 2780 20936
rect 2832 20924 2838 20936
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 2832 20896 4077 20924
rect 2832 20884 2838 20896
rect 4065 20893 4077 20896
rect 4111 20893 4123 20927
rect 6546 20924 6552 20936
rect 6507 20896 6552 20924
rect 4065 20887 4123 20893
rect 6546 20884 6552 20896
rect 6604 20884 6610 20936
rect 9585 20927 9643 20933
rect 9585 20924 9597 20927
rect 9048 20896 9597 20924
rect 3418 20856 3424 20868
rect 3379 20828 3424 20856
rect 3418 20816 3424 20828
rect 3476 20856 3482 20868
rect 4246 20856 4252 20868
rect 3476 20828 4252 20856
rect 3476 20816 3482 20828
rect 4246 20816 4252 20828
rect 4304 20816 4310 20868
rect 5994 20856 6000 20868
rect 5566 20828 6000 20856
rect 5994 20816 6000 20828
rect 6052 20816 6058 20868
rect 6454 20816 6460 20868
rect 6512 20856 6518 20868
rect 6825 20859 6883 20865
rect 6825 20856 6837 20859
rect 6512 20828 6837 20856
rect 6512 20816 6518 20828
rect 6825 20825 6837 20828
rect 6871 20825 6883 20859
rect 8202 20856 8208 20868
rect 8050 20828 8208 20856
rect 6825 20819 6883 20825
rect 8202 20816 8208 20828
rect 8260 20816 8266 20868
rect 8573 20859 8631 20865
rect 8573 20825 8585 20859
rect 8619 20856 8631 20859
rect 8662 20856 8668 20868
rect 8619 20828 8668 20856
rect 8619 20825 8631 20828
rect 8573 20819 8631 20825
rect 8662 20816 8668 20828
rect 8720 20816 8726 20868
rect 9048 20856 9076 20896
rect 9585 20893 9597 20896
rect 9631 20893 9643 20927
rect 9585 20887 9643 20893
rect 9950 20884 9956 20936
rect 10008 20924 10014 20936
rect 10888 20933 10916 20964
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12492 20964 12909 20992
rect 12492 20952 12498 20964
rect 12897 20961 12909 20964
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 12986 20952 12992 21004
rect 13044 20992 13050 21004
rect 13354 20992 13360 21004
rect 13044 20964 13360 20992
rect 13044 20952 13050 20964
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 15304 20992 15332 21032
rect 15378 21020 15384 21072
rect 15436 21060 15442 21072
rect 16206 21060 16212 21072
rect 15436 21032 16212 21060
rect 15436 21020 15442 21032
rect 16206 21020 16212 21032
rect 16264 21020 16270 21072
rect 16482 20992 16488 21004
rect 15304 20964 16488 20992
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 18064 20964 22094 20992
rect 10413 20927 10471 20933
rect 10413 20924 10425 20927
rect 10008 20896 10425 20924
rect 10008 20884 10014 20896
rect 10413 20893 10425 20896
rect 10459 20893 10471 20927
rect 10413 20887 10471 20893
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20893 10931 20927
rect 10873 20887 10931 20893
rect 8772 20828 9076 20856
rect 1854 20748 1860 20800
rect 1912 20788 1918 20800
rect 8772 20788 8800 20828
rect 9398 20816 9404 20868
rect 9456 20856 9462 20868
rect 10888 20856 10916 20887
rect 11238 20884 11244 20936
rect 11296 20924 11302 20936
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 11296 20896 11529 20924
rect 11296 20884 11302 20896
rect 11517 20893 11529 20896
rect 11563 20893 11575 20927
rect 11517 20887 11575 20893
rect 12161 20927 12219 20933
rect 12161 20893 12173 20927
rect 12207 20893 12219 20927
rect 12161 20887 12219 20893
rect 9456 20828 10916 20856
rect 9456 20816 9462 20828
rect 10962 20816 10968 20868
rect 11020 20856 11026 20868
rect 12176 20856 12204 20887
rect 13630 20884 13636 20936
rect 13688 20924 13694 20936
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 13688 20896 14473 20924
rect 13688 20884 13694 20896
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 14550 20884 14556 20936
rect 14608 20924 14614 20936
rect 16390 20924 16396 20936
rect 14608 20896 14653 20924
rect 16351 20896 16396 20924
rect 14608 20884 14614 20896
rect 16390 20884 16396 20896
rect 16448 20884 16454 20936
rect 16850 20924 16856 20936
rect 16811 20896 16856 20924
rect 16850 20884 16856 20896
rect 16908 20924 16914 20936
rect 17497 20927 17555 20933
rect 17497 20924 17509 20927
rect 16908 20896 17509 20924
rect 16908 20884 16914 20896
rect 17497 20893 17509 20896
rect 17543 20893 17555 20927
rect 17497 20887 17555 20893
rect 11020 20828 12204 20856
rect 12989 20859 13047 20865
rect 11020 20816 11026 20828
rect 12989 20825 13001 20859
rect 13035 20856 13047 20859
rect 13078 20856 13084 20868
rect 13035 20828 13084 20856
rect 13035 20825 13047 20828
rect 12989 20819 13047 20825
rect 13078 20816 13084 20828
rect 13136 20816 13142 20868
rect 15013 20859 15071 20865
rect 15013 20825 15025 20859
rect 15059 20856 15071 20859
rect 15378 20856 15384 20868
rect 15059 20828 15384 20856
rect 15059 20825 15071 20828
rect 15013 20819 15071 20825
rect 1912 20760 8800 20788
rect 1912 20748 1918 20760
rect 8938 20748 8944 20800
rect 8996 20788 9002 20800
rect 11238 20788 11244 20800
rect 8996 20760 11244 20788
rect 8996 20748 9002 20760
rect 11238 20748 11244 20760
rect 11296 20748 11302 20800
rect 11609 20791 11667 20797
rect 11609 20757 11621 20791
rect 11655 20788 11667 20791
rect 11882 20788 11888 20800
rect 11655 20760 11888 20788
rect 11655 20757 11667 20760
rect 11609 20751 11667 20757
rect 11882 20748 11888 20760
rect 11940 20748 11946 20800
rect 12710 20748 12716 20800
rect 12768 20788 12774 20800
rect 15028 20788 15056 20819
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 15562 20856 15568 20868
rect 15523 20828 15568 20856
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 15657 20859 15715 20865
rect 15657 20825 15669 20859
rect 15703 20825 15715 20859
rect 16408 20856 16436 20884
rect 18064 20865 18092 20964
rect 18049 20859 18107 20865
rect 18049 20856 18061 20859
rect 16408 20828 18061 20856
rect 15657 20819 15715 20825
rect 18049 20825 18061 20828
rect 18095 20825 18107 20859
rect 18049 20819 18107 20825
rect 12768 20760 15056 20788
rect 15672 20788 15700 20819
rect 19242 20816 19248 20868
rect 19300 20856 19306 20868
rect 19429 20859 19487 20865
rect 19429 20856 19441 20859
rect 19300 20828 19441 20856
rect 19300 20816 19306 20828
rect 19429 20825 19441 20828
rect 19475 20825 19487 20859
rect 19429 20819 19487 20825
rect 19981 20859 20039 20865
rect 19981 20825 19993 20859
rect 20027 20825 20039 20859
rect 19981 20819 20039 20825
rect 20073 20859 20131 20865
rect 20073 20825 20085 20859
rect 20119 20856 20131 20859
rect 21818 20856 21824 20868
rect 20119 20828 21824 20856
rect 20119 20825 20131 20828
rect 20073 20819 20131 20825
rect 16298 20788 16304 20800
rect 15672 20760 16304 20788
rect 12768 20748 12774 20760
rect 16298 20748 16304 20760
rect 16356 20748 16362 20800
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 19996 20788 20024 20819
rect 21818 20816 21824 20828
rect 21876 20816 21882 20868
rect 19392 20760 20024 20788
rect 22066 20788 22094 20964
rect 36170 20788 36176 20800
rect 22066 20760 36176 20788
rect 19392 20748 19398 20760
rect 36170 20748 36176 20760
rect 36228 20748 36234 20800
rect 1104 20698 36892 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 36892 20698
rect 1104 20624 36892 20646
rect 2774 20584 2780 20596
rect 1688 20556 2780 20584
rect 1688 20457 1716 20556
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 3418 20584 3424 20596
rect 3379 20556 3424 20584
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 10226 20584 10232 20596
rect 4080 20556 10232 20584
rect 4080 20516 4108 20556
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 10410 20584 10416 20596
rect 10371 20556 10416 20584
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 11057 20587 11115 20593
rect 11057 20553 11069 20587
rect 11103 20584 11115 20587
rect 13722 20584 13728 20596
rect 11103 20556 13728 20584
rect 11103 20553 11115 20556
rect 11057 20547 11115 20553
rect 13722 20544 13728 20556
rect 13780 20544 13786 20596
rect 14918 20584 14924 20596
rect 14384 20556 14924 20584
rect 4246 20516 4252 20528
rect 3174 20488 4108 20516
rect 4207 20488 4252 20516
rect 4246 20476 4252 20488
rect 4304 20516 4310 20528
rect 5350 20516 5356 20528
rect 4304 20488 5356 20516
rect 4304 20476 4310 20488
rect 5350 20476 5356 20488
rect 5408 20476 5414 20528
rect 5534 20476 5540 20528
rect 5592 20516 5598 20528
rect 6454 20516 6460 20528
rect 5592 20488 6460 20516
rect 5592 20476 5598 20488
rect 6454 20476 6460 20488
rect 6512 20476 6518 20528
rect 6822 20516 6828 20528
rect 6783 20488 6828 20516
rect 6822 20476 6828 20488
rect 6880 20476 6886 20528
rect 6914 20476 6920 20528
rect 6972 20516 6978 20528
rect 7466 20516 7472 20528
rect 6972 20488 7472 20516
rect 6972 20476 6978 20488
rect 7466 20476 7472 20488
rect 7524 20476 7530 20528
rect 10778 20516 10784 20528
rect 8786 20488 10784 20516
rect 10778 20476 10784 20488
rect 10836 20476 10842 20528
rect 12434 20476 12440 20528
rect 12492 20516 12498 20528
rect 12805 20519 12863 20525
rect 12805 20516 12817 20519
rect 12492 20488 12817 20516
rect 12492 20476 12498 20488
rect 12805 20485 12817 20488
rect 12851 20485 12863 20519
rect 12805 20479 12863 20485
rect 12894 20476 12900 20528
rect 12952 20516 12958 20528
rect 13449 20519 13507 20525
rect 12952 20488 12997 20516
rect 12952 20476 12958 20488
rect 13449 20485 13461 20519
rect 13495 20516 13507 20519
rect 14384 20516 14412 20556
rect 14918 20544 14924 20556
rect 14976 20544 14982 20596
rect 15194 20584 15200 20596
rect 15155 20556 15200 20584
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 15654 20544 15660 20596
rect 15712 20584 15718 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 15712 20556 16865 20584
rect 15712 20544 15718 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 20349 20587 20407 20593
rect 20349 20553 20361 20587
rect 20395 20584 20407 20587
rect 23290 20584 23296 20596
rect 20395 20556 23296 20584
rect 20395 20553 20407 20556
rect 20349 20547 20407 20553
rect 13495 20488 14412 20516
rect 14461 20519 14519 20525
rect 13495 20485 13507 20488
rect 13449 20479 13507 20485
rect 14461 20485 14473 20519
rect 14507 20516 14519 20519
rect 15102 20516 15108 20528
rect 14507 20488 15108 20516
rect 14507 20485 14519 20488
rect 14461 20479 14519 20485
rect 15102 20476 15108 20488
rect 15160 20476 15166 20528
rect 16758 20516 16764 20528
rect 15304 20488 16764 20516
rect 15304 20460 15332 20488
rect 16758 20476 16764 20488
rect 16816 20476 16822 20528
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9309 20451 9367 20457
rect 9309 20448 9321 20451
rect 9180 20420 9321 20448
rect 9180 20408 9186 20420
rect 9309 20417 9321 20420
rect 9355 20417 9367 20451
rect 9309 20411 9367 20417
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 10042 20448 10048 20460
rect 9824 20420 10048 20448
rect 9824 20408 9830 20420
rect 10042 20408 10048 20420
rect 10100 20408 10106 20460
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10376 20420 10517 20448
rect 10376 20408 10382 20420
rect 10505 20417 10517 20420
rect 10551 20448 10563 20451
rect 10594 20448 10600 20460
rect 10551 20420 10600 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 10686 20408 10692 20460
rect 10744 20448 10750 20460
rect 10965 20451 11023 20457
rect 10965 20448 10977 20451
rect 10744 20420 10977 20448
rect 10744 20408 10750 20420
rect 10965 20417 10977 20420
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 12069 20451 12127 20457
rect 12069 20417 12081 20451
rect 12115 20448 12127 20451
rect 12342 20448 12348 20460
rect 12115 20420 12348 20448
rect 12115 20417 12127 20420
rect 12069 20411 12127 20417
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 15286 20448 15292 20460
rect 15199 20420 15292 20448
rect 15286 20408 15292 20420
rect 15344 20408 15350 20460
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20448 16267 20451
rect 16574 20448 16580 20460
rect 16255 20420 16580 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 16868 20448 16896 20547
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 35989 20587 36047 20593
rect 35989 20553 36001 20587
rect 36035 20584 36047 20587
rect 36078 20584 36084 20596
rect 36035 20556 36084 20584
rect 36035 20553 36047 20556
rect 35989 20547 36047 20553
rect 36078 20544 36084 20556
rect 36136 20544 36142 20596
rect 17405 20451 17463 20457
rect 17405 20448 17417 20451
rect 16868 20420 17417 20448
rect 17405 20417 17417 20420
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20448 20223 20451
rect 20254 20448 20260 20460
rect 20211 20420 20260 20448
rect 20211 20417 20223 20420
rect 20165 20411 20223 20417
rect 20254 20408 20260 20420
rect 20312 20448 20318 20460
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 20312 20420 20821 20448
rect 20312 20408 20318 20420
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 35805 20451 35863 20457
rect 35805 20448 35817 20451
rect 20809 20411 20867 20417
rect 35268 20420 35817 20448
rect 1949 20383 2007 20389
rect 1949 20349 1961 20383
rect 1995 20380 2007 20383
rect 2958 20380 2964 20392
rect 1995 20352 2964 20380
rect 1995 20349 2007 20352
rect 1949 20343 2007 20349
rect 2958 20340 2964 20352
rect 3016 20380 3022 20392
rect 3326 20380 3332 20392
rect 3016 20352 3332 20380
rect 3016 20340 3022 20352
rect 3326 20340 3332 20352
rect 3384 20340 3390 20392
rect 5902 20380 5908 20392
rect 5863 20352 5908 20380
rect 5902 20340 5908 20352
rect 5960 20380 5966 20392
rect 6546 20380 6552 20392
rect 5960 20352 6552 20380
rect 5960 20340 5966 20352
rect 6546 20340 6552 20352
rect 6604 20380 6610 20392
rect 7190 20380 7196 20392
rect 6604 20352 7196 20380
rect 6604 20340 6610 20352
rect 7190 20340 7196 20352
rect 7248 20380 7254 20392
rect 7285 20383 7343 20389
rect 7285 20380 7297 20383
rect 7248 20352 7297 20380
rect 7248 20340 7254 20352
rect 7285 20349 7297 20352
rect 7331 20349 7343 20383
rect 7285 20343 7343 20349
rect 7561 20383 7619 20389
rect 7561 20349 7573 20383
rect 7607 20380 7619 20383
rect 8754 20380 8760 20392
rect 7607 20352 8760 20380
rect 7607 20349 7619 20352
rect 7561 20343 7619 20349
rect 8754 20340 8760 20352
rect 8812 20340 8818 20392
rect 8846 20340 8852 20392
rect 8904 20380 8910 20392
rect 11790 20380 11796 20392
rect 8904 20352 11796 20380
rect 8904 20340 8910 20352
rect 11790 20340 11796 20352
rect 11848 20340 11854 20392
rect 12526 20380 12532 20392
rect 12406 20352 12532 20380
rect 12406 20312 12434 20352
rect 12526 20340 12532 20352
rect 12584 20340 12590 20392
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 14553 20383 14611 20389
rect 14553 20380 14565 20383
rect 13504 20352 14565 20380
rect 13504 20340 13510 20352
rect 14553 20349 14565 20352
rect 14599 20349 14611 20383
rect 19153 20383 19211 20389
rect 19153 20380 19165 20383
rect 14553 20343 14611 20349
rect 14660 20352 19165 20380
rect 10060 20284 12434 20312
rect 14001 20315 14059 20321
rect 10060 20256 10088 20284
rect 14001 20281 14013 20315
rect 14047 20312 14059 20315
rect 14274 20312 14280 20324
rect 14047 20284 14280 20312
rect 14047 20281 14059 20284
rect 14001 20275 14059 20281
rect 14274 20272 14280 20284
rect 14332 20272 14338 20324
rect 6730 20204 6736 20256
rect 6788 20244 6794 20256
rect 9398 20244 9404 20256
rect 6788 20216 9404 20244
rect 6788 20204 6794 20216
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 9861 20247 9919 20253
rect 9861 20213 9873 20247
rect 9907 20244 9919 20247
rect 10042 20244 10048 20256
rect 9907 20216 10048 20244
rect 9907 20213 9919 20216
rect 9861 20207 9919 20213
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 12161 20247 12219 20253
rect 12161 20213 12173 20247
rect 12207 20244 12219 20247
rect 12618 20244 12624 20256
rect 12207 20216 12624 20244
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 12618 20204 12624 20216
rect 12676 20204 12682 20256
rect 12710 20204 12716 20256
rect 12768 20244 12774 20256
rect 14660 20244 14688 20352
rect 19153 20349 19165 20352
rect 19199 20349 19211 20383
rect 19153 20343 19211 20349
rect 16022 20312 16028 20324
rect 15983 20284 16028 20312
rect 16022 20272 16028 20284
rect 16080 20272 16086 20324
rect 17497 20315 17555 20321
rect 17497 20281 17509 20315
rect 17543 20312 17555 20315
rect 19610 20312 19616 20324
rect 17543 20284 19616 20312
rect 17543 20281 17555 20284
rect 17497 20275 17555 20281
rect 19610 20272 19616 20284
rect 19668 20272 19674 20324
rect 12768 20216 14688 20244
rect 12768 20204 12774 20216
rect 14918 20204 14924 20256
rect 14976 20244 14982 20256
rect 17218 20244 17224 20256
rect 14976 20216 17224 20244
rect 14976 20204 14982 20216
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 18141 20247 18199 20253
rect 18141 20213 18153 20247
rect 18187 20244 18199 20247
rect 18414 20244 18420 20256
rect 18187 20216 18420 20244
rect 18187 20213 18199 20216
rect 18141 20207 18199 20213
rect 18414 20204 18420 20216
rect 18472 20244 18478 20256
rect 18601 20247 18659 20253
rect 18601 20244 18613 20247
rect 18472 20216 18613 20244
rect 18472 20204 18478 20216
rect 18601 20213 18613 20216
rect 18647 20213 18659 20247
rect 18601 20207 18659 20213
rect 34514 20204 34520 20256
rect 34572 20244 34578 20256
rect 35268 20253 35296 20420
rect 35805 20417 35817 20420
rect 35851 20417 35863 20451
rect 35805 20411 35863 20417
rect 35253 20247 35311 20253
rect 35253 20244 35265 20247
rect 34572 20216 35265 20244
rect 34572 20204 34578 20216
rect 35253 20213 35265 20216
rect 35299 20213 35311 20247
rect 35253 20207 35311 20213
rect 1104 20154 36892 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 36892 20154
rect 1104 20080 36892 20102
rect 1673 20043 1731 20049
rect 1673 20009 1685 20043
rect 1719 20040 1731 20043
rect 1762 20040 1768 20052
rect 1719 20012 1768 20040
rect 1719 20009 1731 20012
rect 1673 20003 1731 20009
rect 1762 20000 1768 20012
rect 1820 20040 1826 20052
rect 2590 20040 2596 20052
rect 1820 20012 2596 20040
rect 1820 20000 1826 20012
rect 2590 20000 2596 20012
rect 2648 20000 2654 20052
rect 3510 20000 3516 20052
rect 3568 20040 3574 20052
rect 5997 20043 6055 20049
rect 3568 20012 5948 20040
rect 3568 20000 3574 20012
rect 5920 19972 5948 20012
rect 5997 20009 6009 20043
rect 6043 20040 6055 20043
rect 6822 20040 6828 20052
rect 6043 20012 6828 20040
rect 6043 20009 6055 20012
rect 5997 20003 6055 20009
rect 6822 20000 6828 20012
rect 6880 20040 6886 20052
rect 7558 20040 7564 20052
rect 6880 20012 7564 20040
rect 6880 20000 6886 20012
rect 7558 20000 7564 20012
rect 7616 20000 7622 20052
rect 7650 20000 7656 20052
rect 7708 20040 7714 20052
rect 7708 20012 8432 20040
rect 7708 20000 7714 20012
rect 8404 19972 8432 20012
rect 8478 20000 8484 20052
rect 8536 20040 8542 20052
rect 8662 20040 8668 20052
rect 8536 20012 8668 20040
rect 8536 20000 8542 20012
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 9858 20040 9864 20052
rect 9819 20012 9864 20040
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10192 20012 13768 20040
rect 10192 20000 10198 20012
rect 9030 19972 9036 19984
rect 5920 19944 6868 19972
rect 8404 19944 9036 19972
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 3421 19907 3479 19913
rect 3421 19904 3433 19907
rect 2832 19876 3433 19904
rect 2832 19864 2838 19876
rect 3421 19873 3433 19876
rect 3467 19904 3479 19907
rect 4062 19904 4068 19916
rect 3467 19876 4068 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 4062 19864 4068 19876
rect 4120 19904 4126 19916
rect 4249 19907 4307 19913
rect 4249 19904 4261 19907
rect 4120 19876 4261 19904
rect 4120 19864 4126 19876
rect 4249 19873 4261 19876
rect 4295 19873 4307 19907
rect 4249 19867 4307 19873
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 4890 19904 4896 19916
rect 4571 19876 4896 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 5902 19864 5908 19916
rect 5960 19904 5966 19916
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 5960 19876 6745 19904
rect 5960 19864 5966 19876
rect 6733 19873 6745 19876
rect 6779 19873 6791 19907
rect 6840 19904 6868 19944
rect 9030 19932 9036 19944
rect 9088 19932 9094 19984
rect 9214 19932 9220 19984
rect 9272 19972 9278 19984
rect 10505 19975 10563 19981
rect 10505 19972 10517 19975
rect 9272 19944 10517 19972
rect 9272 19932 9278 19944
rect 10505 19941 10517 19944
rect 10551 19941 10563 19975
rect 11974 19972 11980 19984
rect 10505 19935 10563 19941
rect 11532 19944 11980 19972
rect 7742 19904 7748 19916
rect 6840 19876 7748 19904
rect 6733 19867 6791 19873
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 8481 19907 8539 19913
rect 8481 19873 8493 19907
rect 8527 19904 8539 19907
rect 11422 19904 11428 19916
rect 8527 19876 11428 19904
rect 8527 19873 8539 19876
rect 8481 19867 8539 19873
rect 11422 19864 11428 19876
rect 11480 19864 11486 19916
rect 9122 19796 9128 19848
rect 9180 19836 9186 19848
rect 9309 19839 9367 19845
rect 9309 19836 9321 19839
rect 9180 19808 9321 19836
rect 9180 19796 9186 19808
rect 9309 19805 9321 19808
rect 9355 19836 9367 19839
rect 9950 19836 9956 19848
rect 9355 19808 9674 19836
rect 9911 19808 9956 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 2682 19728 2688 19780
rect 2740 19728 2746 19780
rect 3145 19771 3203 19777
rect 3145 19737 3157 19771
rect 3191 19737 3203 19771
rect 5750 19740 6684 19768
rect 3145 19731 3203 19737
rect 3160 19700 3188 19731
rect 6454 19700 6460 19712
rect 3160 19672 6460 19700
rect 6454 19660 6460 19672
rect 6512 19660 6518 19712
rect 6656 19700 6684 19740
rect 6730 19728 6736 19780
rect 6788 19768 6794 19780
rect 7009 19771 7067 19777
rect 7009 19768 7021 19771
rect 6788 19740 7021 19768
rect 6788 19728 6794 19740
rect 7009 19737 7021 19740
rect 7055 19737 7067 19771
rect 9217 19771 9275 19777
rect 9217 19768 9229 19771
rect 8234 19740 9229 19768
rect 7009 19731 7067 19737
rect 9217 19737 9229 19740
rect 9263 19737 9275 19771
rect 9646 19768 9674 19808
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 10870 19836 10876 19848
rect 10643 19808 10876 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 10410 19768 10416 19780
rect 9646 19740 10416 19768
rect 9217 19731 9275 19737
rect 10410 19728 10416 19740
rect 10468 19768 10474 19780
rect 10612 19768 10640 19799
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19836 11115 19839
rect 11532 19836 11560 19944
rect 11974 19932 11980 19944
rect 12032 19932 12038 19984
rect 12345 19975 12403 19981
rect 12345 19941 12357 19975
rect 12391 19972 12403 19975
rect 13740 19972 13768 20012
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14369 20043 14427 20049
rect 14369 20040 14381 20043
rect 13872 20012 14381 20040
rect 13872 20000 13878 20012
rect 14369 20009 14381 20012
rect 14415 20009 14427 20043
rect 15102 20040 15108 20052
rect 15063 20012 15108 20040
rect 14369 20003 14427 20009
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 16850 20040 16856 20052
rect 15212 20012 16856 20040
rect 15212 19972 15240 20012
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 17126 20000 17132 20052
rect 17184 20040 17190 20052
rect 17497 20043 17555 20049
rect 17497 20040 17509 20043
rect 17184 20012 17509 20040
rect 17184 20000 17190 20012
rect 17497 20009 17509 20012
rect 17543 20009 17555 20043
rect 17497 20003 17555 20009
rect 20254 20000 20260 20052
rect 20312 20040 20318 20052
rect 36630 20040 36636 20052
rect 20312 20012 36636 20040
rect 20312 20000 20318 20012
rect 36630 20000 36636 20012
rect 36688 20000 36694 20052
rect 17310 19972 17316 19984
rect 12391 19944 13676 19972
rect 13740 19944 15240 19972
rect 12391 19941 12403 19944
rect 12345 19935 12403 19941
rect 11790 19904 11796 19916
rect 11751 19876 11796 19904
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 12158 19864 12164 19916
rect 12216 19904 12222 19916
rect 12897 19907 12955 19913
rect 12897 19904 12909 19907
rect 12216 19876 12909 19904
rect 12216 19864 12222 19876
rect 12897 19873 12909 19876
rect 12943 19873 12955 19907
rect 12897 19867 12955 19873
rect 13446 19864 13452 19916
rect 13504 19904 13510 19916
rect 13541 19907 13599 19913
rect 13541 19904 13553 19907
rect 13504 19876 13553 19904
rect 13504 19864 13510 19876
rect 13541 19873 13553 19876
rect 13587 19873 13599 19907
rect 13648 19904 13676 19944
rect 14274 19904 14280 19916
rect 13648 19876 14280 19904
rect 13541 19867 13599 19873
rect 14274 19864 14280 19876
rect 14332 19864 14338 19916
rect 14458 19836 14464 19848
rect 11103 19808 11560 19836
rect 14419 19808 14464 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 10468 19740 10640 19768
rect 10468 19728 10474 19740
rect 8294 19700 8300 19712
rect 6656 19672 8300 19700
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 9030 19660 9036 19712
rect 9088 19700 9094 19712
rect 11072 19700 11100 19799
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 15212 19845 15240 19944
rect 15764 19944 17316 19972
rect 15197 19839 15255 19845
rect 15197 19805 15209 19839
rect 15243 19805 15255 19839
rect 15197 19799 15255 19805
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 11940 19740 11985 19768
rect 11940 19728 11946 19740
rect 12066 19728 12072 19780
rect 12124 19768 12130 19780
rect 13446 19768 13452 19780
rect 12124 19740 13308 19768
rect 13407 19740 13452 19768
rect 12124 19728 12130 19740
rect 9088 19672 11100 19700
rect 11149 19703 11207 19709
rect 9088 19660 9094 19672
rect 11149 19669 11161 19703
rect 11195 19700 11207 19703
rect 13078 19700 13084 19712
rect 11195 19672 13084 19700
rect 11195 19669 11207 19672
rect 11149 19663 11207 19669
rect 13078 19660 13084 19672
rect 13136 19660 13142 19712
rect 13280 19700 13308 19740
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 13722 19728 13728 19780
rect 13780 19768 13786 19780
rect 15764 19768 15792 19944
rect 17310 19932 17316 19944
rect 17368 19972 17374 19984
rect 18785 19975 18843 19981
rect 18785 19972 18797 19975
rect 17368 19944 18797 19972
rect 17368 19932 17374 19944
rect 18785 19941 18797 19944
rect 18831 19972 18843 19975
rect 19058 19972 19064 19984
rect 18831 19944 19064 19972
rect 18831 19941 18843 19944
rect 18785 19935 18843 19941
rect 19058 19932 19064 19944
rect 19116 19932 19122 19984
rect 19426 19932 19432 19984
rect 19484 19972 19490 19984
rect 19484 19944 19564 19972
rect 19484 19932 19490 19944
rect 19536 19913 19564 19944
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 20438 19904 20444 19916
rect 19567 19876 20444 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19836 15899 19839
rect 16945 19839 17003 19845
rect 15887 19808 16436 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 13780 19740 15792 19768
rect 13780 19728 13786 19740
rect 14366 19700 14372 19712
rect 13280 19672 14372 19700
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 15194 19660 15200 19712
rect 15252 19700 15258 19712
rect 16408 19709 16436 19808
rect 16945 19805 16957 19839
rect 16991 19836 17003 19839
rect 17589 19839 17647 19845
rect 17589 19836 17601 19839
rect 16991 19808 17601 19836
rect 16991 19805 17003 19808
rect 16945 19799 17003 19805
rect 17589 19805 17601 19808
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19836 18291 19839
rect 18414 19836 18420 19848
rect 18279 19808 18420 19836
rect 18279 19805 18291 19808
rect 18233 19799 18291 19805
rect 17604 19768 17632 19799
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 22462 19836 22468 19848
rect 22423 19808 22468 19836
rect 22462 19796 22468 19808
rect 22520 19836 22526 19848
rect 22922 19836 22928 19848
rect 22520 19808 22928 19836
rect 22520 19796 22526 19808
rect 22922 19796 22928 19808
rect 22980 19796 22986 19848
rect 18598 19768 18604 19780
rect 17604 19740 18604 19768
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 19610 19728 19616 19780
rect 19668 19768 19674 19780
rect 20162 19768 20168 19780
rect 19668 19740 19713 19768
rect 20075 19740 20168 19768
rect 19668 19728 19674 19740
rect 20162 19728 20168 19740
rect 20220 19768 20226 19780
rect 20530 19768 20536 19780
rect 20220 19740 20536 19768
rect 20220 19728 20226 19740
rect 20530 19728 20536 19740
rect 20588 19728 20594 19780
rect 15749 19703 15807 19709
rect 15749 19700 15761 19703
rect 15252 19672 15761 19700
rect 15252 19660 15258 19672
rect 15749 19669 15761 19672
rect 15795 19669 15807 19703
rect 15749 19663 15807 19669
rect 16393 19703 16451 19709
rect 16393 19669 16405 19703
rect 16439 19700 16451 19703
rect 16574 19700 16580 19712
rect 16439 19672 16580 19700
rect 16439 19669 16451 19672
rect 16393 19663 16451 19669
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 18138 19700 18144 19712
rect 18099 19672 18144 19700
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 22186 19660 22192 19712
rect 22244 19700 22250 19712
rect 22373 19703 22431 19709
rect 22373 19700 22385 19703
rect 22244 19672 22385 19700
rect 22244 19660 22250 19672
rect 22373 19669 22385 19672
rect 22419 19669 22431 19703
rect 22373 19663 22431 19669
rect 1104 19610 36892 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 36892 19610
rect 1104 19536 36892 19558
rect 5534 19496 5540 19508
rect 3620 19468 5540 19496
rect 3510 19428 3516 19440
rect 3082 19400 3516 19428
rect 3510 19388 3516 19400
rect 3568 19388 3574 19440
rect 3620 19437 3648 19468
rect 5534 19456 5540 19468
rect 5592 19456 5598 19508
rect 5810 19456 5816 19508
rect 5868 19496 5874 19508
rect 5997 19499 6055 19505
rect 5997 19496 6009 19499
rect 5868 19468 6009 19496
rect 5868 19456 5874 19468
rect 5997 19465 6009 19468
rect 6043 19465 6055 19499
rect 5997 19459 6055 19465
rect 6454 19456 6460 19508
rect 6512 19496 6518 19508
rect 7650 19496 7656 19508
rect 6512 19468 7656 19496
rect 6512 19456 6518 19468
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 8570 19496 8576 19508
rect 7760 19468 8576 19496
rect 3605 19431 3663 19437
rect 3605 19397 3617 19431
rect 3651 19397 3663 19431
rect 7466 19428 7472 19440
rect 5750 19400 7472 19428
rect 3605 19391 3663 19397
rect 7466 19388 7472 19400
rect 7524 19388 7530 19440
rect 7760 19437 7788 19468
rect 8570 19456 8576 19468
rect 8628 19496 8634 19508
rect 8754 19496 8760 19508
rect 8628 19468 8760 19496
rect 8628 19456 8634 19468
rect 8754 19456 8760 19468
rect 8812 19456 8818 19508
rect 11885 19499 11943 19505
rect 11885 19465 11897 19499
rect 11931 19496 11943 19499
rect 11931 19468 13400 19496
rect 11931 19465 11943 19468
rect 11885 19459 11943 19465
rect 7745 19431 7803 19437
rect 7745 19397 7757 19431
rect 7791 19397 7803 19431
rect 9582 19428 9588 19440
rect 8970 19400 9588 19428
rect 7745 19391 7803 19397
rect 9582 19388 9588 19400
rect 9640 19388 9646 19440
rect 12618 19428 12624 19440
rect 10336 19400 12388 19428
rect 12579 19400 12624 19428
rect 1578 19360 1584 19372
rect 1539 19332 1584 19360
rect 1578 19320 1584 19332
rect 1636 19320 1642 19372
rect 4062 19320 4068 19372
rect 4120 19360 4126 19372
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 4120 19332 4261 19360
rect 4120 19320 4126 19332
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 6914 19360 6920 19372
rect 6875 19332 6920 19360
rect 4249 19323 4307 19329
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19360 7067 19363
rect 7098 19360 7104 19372
rect 7055 19332 7104 19360
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 9456 19332 9505 19360
rect 9456 19320 9462 19332
rect 9493 19329 9505 19332
rect 9539 19360 9551 19363
rect 10336 19360 10364 19400
rect 9539 19332 10364 19360
rect 9539 19329 9551 19332
rect 9493 19323 9551 19329
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 10505 19363 10563 19369
rect 10505 19360 10517 19363
rect 10468 19332 10517 19360
rect 10468 19320 10474 19332
rect 10505 19329 10517 19332
rect 10551 19329 10563 19363
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10505 19323 10563 19329
rect 10612 19332 10977 19360
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19292 1915 19295
rect 1946 19292 1952 19304
rect 1903 19264 1952 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 4522 19292 4528 19304
rect 4483 19264 4528 19292
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 5258 19252 5264 19304
rect 5316 19292 5322 19304
rect 7190 19292 7196 19304
rect 5316 19264 7196 19292
rect 5316 19252 5322 19264
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 7282 19252 7288 19304
rect 7340 19292 7346 19304
rect 7469 19295 7527 19301
rect 7469 19292 7481 19295
rect 7340 19264 7481 19292
rect 7340 19252 7346 19264
rect 7469 19261 7481 19264
rect 7515 19261 7527 19295
rect 10612 19292 10640 19332
rect 10965 19329 10977 19332
rect 11011 19360 11023 19363
rect 11011 19332 11376 19360
rect 11011 19329 11023 19332
rect 10965 19323 11023 19329
rect 7469 19255 7527 19261
rect 7576 19264 10640 19292
rect 11348 19292 11376 19332
rect 11422 19320 11428 19372
rect 11480 19360 11486 19372
rect 11793 19363 11851 19369
rect 11793 19360 11805 19363
rect 11480 19332 11805 19360
rect 11480 19320 11486 19332
rect 11793 19329 11805 19332
rect 11839 19329 11851 19363
rect 12066 19360 12072 19372
rect 11793 19323 11851 19329
rect 11900 19332 12072 19360
rect 11900 19292 11928 19332
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 11348 19264 11928 19292
rect 5534 19184 5540 19236
rect 5592 19224 5598 19236
rect 7006 19224 7012 19236
rect 5592 19196 7012 19224
rect 5592 19184 5598 19196
rect 7006 19184 7012 19196
rect 7064 19184 7070 19236
rect 7098 19184 7104 19236
rect 7156 19224 7162 19236
rect 7374 19224 7380 19236
rect 7156 19196 7380 19224
rect 7156 19184 7162 19196
rect 7374 19184 7380 19196
rect 7432 19224 7438 19236
rect 7576 19224 7604 19264
rect 7432 19196 7604 19224
rect 7432 19184 7438 19196
rect 8754 19184 8760 19236
rect 8812 19224 8818 19236
rect 11882 19224 11888 19236
rect 8812 19196 11888 19224
rect 8812 19184 8818 19196
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 12360 19224 12388 19400
rect 12618 19388 12624 19400
rect 12676 19388 12682 19440
rect 13372 19428 13400 19468
rect 13446 19456 13452 19508
rect 13504 19496 13510 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 13504 19468 14933 19496
rect 13504 19456 13510 19468
rect 14921 19465 14933 19468
rect 14967 19465 14979 19499
rect 14921 19459 14979 19465
rect 16114 19456 16120 19508
rect 16172 19496 16178 19508
rect 16209 19499 16267 19505
rect 16209 19496 16221 19499
rect 16172 19468 16221 19496
rect 16172 19456 16178 19468
rect 16209 19465 16221 19468
rect 16255 19465 16267 19499
rect 18509 19499 18567 19505
rect 16209 19459 16267 19465
rect 16316 19468 18276 19496
rect 14826 19428 14832 19440
rect 13372 19400 14832 19428
rect 14826 19388 14832 19400
rect 14884 19388 14890 19440
rect 16316 19428 16344 19468
rect 14936 19400 16344 19428
rect 17037 19431 17095 19437
rect 13538 19320 13544 19372
rect 13596 19360 13602 19372
rect 14277 19363 14335 19369
rect 14277 19360 14289 19363
rect 13596 19332 14289 19360
rect 13596 19320 13602 19332
rect 14277 19329 14289 19332
rect 14323 19329 14335 19363
rect 14277 19323 14335 19329
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19360 14427 19363
rect 14642 19360 14648 19372
rect 14415 19332 14648 19360
rect 14415 19329 14427 19332
rect 14369 19323 14427 19329
rect 14642 19320 14648 19332
rect 14700 19360 14706 19372
rect 14936 19360 14964 19400
rect 17037 19397 17049 19431
rect 17083 19428 17095 19431
rect 18138 19428 18144 19440
rect 17083 19400 18144 19428
rect 17083 19397 17095 19400
rect 17037 19391 17095 19397
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 18248 19428 18276 19468
rect 18509 19465 18521 19499
rect 18555 19496 18567 19499
rect 19334 19496 19340 19508
rect 18555 19468 19340 19496
rect 18555 19465 18567 19468
rect 18509 19459 18567 19465
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 18782 19428 18788 19440
rect 18248 19400 18788 19428
rect 18782 19388 18788 19400
rect 18840 19388 18846 19440
rect 19981 19431 20039 19437
rect 19981 19397 19993 19431
rect 20027 19428 20039 19431
rect 21266 19428 21272 19440
rect 20027 19400 21272 19428
rect 20027 19397 20039 19400
rect 19981 19391 20039 19397
rect 21266 19388 21272 19400
rect 21324 19388 21330 19440
rect 22186 19428 22192 19440
rect 22147 19400 22192 19428
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 14700 19332 14964 19360
rect 14700 19320 14706 19332
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 15657 19363 15715 19369
rect 15068 19332 15113 19360
rect 15068 19320 15074 19332
rect 15657 19329 15669 19363
rect 15703 19360 15715 19363
rect 15930 19360 15936 19372
rect 15703 19332 15936 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 16114 19320 16120 19372
rect 16172 19360 16178 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 16172 19332 16313 19360
rect 16172 19320 16178 19332
rect 16301 19329 16313 19332
rect 16347 19360 16359 19363
rect 16390 19360 16396 19372
rect 16347 19332 16396 19360
rect 16347 19329 16359 19332
rect 16301 19323 16359 19329
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 19058 19360 19064 19372
rect 19019 19332 19064 19360
rect 19058 19320 19064 19332
rect 19116 19320 19122 19372
rect 19153 19363 19211 19369
rect 19153 19329 19165 19363
rect 19199 19360 19211 19363
rect 19702 19360 19708 19372
rect 19199 19332 19708 19360
rect 19199 19329 19211 19332
rect 19153 19323 19211 19329
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 35894 19320 35900 19372
rect 35952 19360 35958 19372
rect 35952 19332 35997 19360
rect 35952 19320 35958 19332
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19292 12587 19295
rect 12710 19292 12716 19304
rect 12575 19264 12716 19292
rect 12575 19261 12587 19264
rect 12529 19255 12587 19261
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 13173 19295 13231 19301
rect 13173 19261 13185 19295
rect 13219 19292 13231 19295
rect 13998 19292 14004 19304
rect 13219 19264 14004 19292
rect 13219 19261 13231 19264
rect 13173 19255 13231 19261
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14918 19292 14924 19304
rect 14792 19264 14924 19292
rect 14792 19252 14798 19264
rect 14918 19252 14924 19264
rect 14976 19292 14982 19304
rect 16942 19292 16948 19304
rect 14976 19264 16436 19292
rect 16903 19264 16948 19292
rect 14976 19252 14982 19264
rect 12434 19224 12440 19236
rect 12360 19196 12440 19224
rect 12434 19184 12440 19196
rect 12492 19224 12498 19236
rect 12802 19224 12808 19236
rect 12492 19196 12808 19224
rect 12492 19184 12498 19196
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 13725 19227 13783 19233
rect 13725 19193 13737 19227
rect 13771 19224 13783 19227
rect 16114 19224 16120 19236
rect 13771 19196 16120 19224
rect 13771 19193 13783 19196
rect 13725 19187 13783 19193
rect 16114 19184 16120 19196
rect 16172 19184 16178 19236
rect 16408 19224 16436 19264
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17221 19295 17279 19301
rect 17221 19261 17233 19295
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 19889 19295 19947 19301
rect 19889 19261 19901 19295
rect 19935 19292 19947 19295
rect 19978 19292 19984 19304
rect 19935 19264 19984 19292
rect 19935 19261 19947 19264
rect 19889 19255 19947 19261
rect 17236 19224 17264 19255
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20165 19295 20223 19301
rect 20165 19261 20177 19295
rect 20211 19261 20223 19295
rect 21082 19292 21088 19304
rect 21043 19264 21088 19292
rect 20165 19255 20223 19261
rect 20180 19224 20208 19255
rect 21082 19252 21088 19264
rect 21140 19252 21146 19304
rect 22094 19292 22100 19304
rect 22055 19264 22100 19292
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 22373 19295 22431 19301
rect 22373 19261 22385 19295
rect 22419 19261 22431 19295
rect 22373 19255 22431 19261
rect 22388 19224 22416 19255
rect 16408 19196 17264 19224
rect 19444 19196 22416 19224
rect 2498 19116 2504 19168
rect 2556 19156 2562 19168
rect 4890 19156 4896 19168
rect 2556 19128 4896 19156
rect 2556 19116 2562 19128
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 9306 19156 9312 19168
rect 5316 19128 9312 19156
rect 5316 19116 5322 19128
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 10410 19156 10416 19168
rect 10371 19128 10416 19156
rect 10410 19116 10416 19128
rect 10468 19116 10474 19168
rect 11057 19159 11115 19165
rect 11057 19125 11069 19159
rect 11103 19156 11115 19159
rect 12066 19156 12072 19168
rect 11103 19128 12072 19156
rect 11103 19125 11115 19128
rect 11057 19119 11115 19125
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 15436 19128 15577 19156
rect 15436 19116 15442 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 15565 19119 15623 19125
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 19444 19156 19472 19196
rect 36078 19156 36084 19168
rect 15896 19128 19472 19156
rect 36039 19128 36084 19156
rect 15896 19116 15902 19128
rect 36078 19116 36084 19128
rect 36136 19116 36142 19168
rect 1104 19066 36892 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 36892 19066
rect 1104 18992 36892 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 1452 18924 1593 18952
rect 1452 18912 1458 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 6086 18952 6092 18964
rect 1581 18915 1639 18921
rect 3252 18924 6092 18952
rect 3053 18819 3111 18825
rect 3053 18785 3065 18819
rect 3099 18816 3111 18819
rect 3252 18816 3280 18924
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 6825 18955 6883 18961
rect 6825 18921 6837 18955
rect 6871 18952 6883 18955
rect 7006 18952 7012 18964
rect 6871 18924 7012 18952
rect 6871 18921 6883 18924
rect 6825 18915 6883 18921
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 7190 18912 7196 18964
rect 7248 18952 7254 18964
rect 9493 18955 9551 18961
rect 9493 18952 9505 18955
rect 7248 18924 9505 18952
rect 7248 18912 7254 18924
rect 9493 18921 9505 18924
rect 9539 18921 9551 18955
rect 14366 18952 14372 18964
rect 14279 18924 14372 18952
rect 9493 18915 9551 18921
rect 14366 18912 14372 18924
rect 14424 18952 14430 18964
rect 15286 18952 15292 18964
rect 14424 18924 15292 18952
rect 14424 18912 14430 18924
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16945 18955 17003 18961
rect 16945 18952 16957 18955
rect 16632 18924 16957 18952
rect 16632 18912 16638 18924
rect 16945 18921 16957 18924
rect 16991 18952 17003 18955
rect 29822 18952 29828 18964
rect 16991 18924 29828 18952
rect 16991 18921 17003 18924
rect 16945 18915 17003 18921
rect 29822 18912 29828 18924
rect 29880 18912 29886 18964
rect 6362 18884 6368 18896
rect 5920 18856 6368 18884
rect 3099 18788 3280 18816
rect 3329 18819 3387 18825
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 4062 18816 4068 18828
rect 3375 18788 4068 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 5166 18816 5172 18828
rect 4540 18788 5172 18816
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18748 4031 18751
rect 4540 18748 4568 18788
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 5626 18776 5632 18828
rect 5684 18816 5690 18828
rect 5721 18819 5779 18825
rect 5721 18816 5733 18819
rect 5684 18788 5733 18816
rect 5684 18776 5690 18788
rect 5721 18785 5733 18788
rect 5767 18816 5779 18819
rect 5920 18816 5948 18856
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 13538 18884 13544 18896
rect 10704 18856 13544 18884
rect 5767 18788 5948 18816
rect 5997 18819 6055 18825
rect 5767 18785 5779 18788
rect 5721 18779 5779 18785
rect 5997 18785 6009 18819
rect 6043 18816 6055 18819
rect 7282 18816 7288 18828
rect 6043 18788 7288 18816
rect 6043 18785 6055 18788
rect 5997 18779 6055 18785
rect 7282 18776 7288 18788
rect 7340 18816 7346 18828
rect 8573 18819 8631 18825
rect 8573 18816 8585 18819
rect 7340 18788 8585 18816
rect 7340 18776 7346 18788
rect 8573 18785 8585 18788
rect 8619 18785 8631 18819
rect 8573 18779 8631 18785
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 10704 18816 10732 18856
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 14148 18856 15792 18884
rect 14148 18844 14154 18856
rect 9916 18788 10732 18816
rect 9916 18776 9922 18788
rect 9582 18748 9588 18760
rect 4019 18720 4568 18748
rect 9543 18720 9588 18748
rect 4019 18717 4031 18720
rect 3973 18711 4031 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 10008 18720 10241 18748
rect 10008 18708 10014 18720
rect 10229 18717 10241 18720
rect 10275 18748 10287 18751
rect 10594 18748 10600 18760
rect 10275 18720 10600 18748
rect 10275 18717 10287 18720
rect 10229 18711 10287 18717
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 10704 18757 10732 18788
rect 11425 18819 11483 18825
rect 11425 18785 11437 18819
rect 11471 18816 11483 18819
rect 11790 18816 11796 18828
rect 11471 18788 11796 18816
rect 11471 18785 11483 18788
rect 11425 18779 11483 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18816 13231 18819
rect 15194 18816 15200 18828
rect 13219 18788 15200 18816
rect 13219 18785 13231 18788
rect 13173 18779 13231 18785
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 15470 18816 15476 18828
rect 15431 18788 15476 18816
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 15764 18748 15792 18856
rect 16482 18844 16488 18896
rect 16540 18884 16546 18896
rect 18233 18887 18291 18893
rect 18233 18884 18245 18887
rect 16540 18856 18245 18884
rect 16540 18844 16546 18856
rect 18233 18853 18245 18856
rect 18279 18884 18291 18887
rect 18279 18856 19564 18884
rect 18279 18853 18291 18856
rect 18233 18847 18291 18853
rect 16393 18819 16451 18825
rect 16393 18785 16405 18819
rect 16439 18816 16451 18819
rect 16942 18816 16948 18828
rect 16439 18788 16948 18816
rect 16439 18785 16451 18788
rect 16393 18779 16451 18785
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 19536 18825 19564 18856
rect 20622 18844 20628 18896
rect 20680 18884 20686 18896
rect 24854 18884 24860 18896
rect 20680 18856 24860 18884
rect 20680 18844 20686 18856
rect 24854 18844 24860 18856
rect 24912 18844 24918 18896
rect 19521 18819 19579 18825
rect 19521 18785 19533 18819
rect 19567 18816 19579 18819
rect 20162 18816 20168 18828
rect 19567 18788 20168 18816
rect 19567 18785 19579 18788
rect 19521 18779 19579 18785
rect 20162 18776 20168 18788
rect 20220 18776 20226 18828
rect 21818 18816 21824 18828
rect 21779 18788 21824 18816
rect 21818 18776 21824 18788
rect 21876 18776 21882 18828
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 15764 18720 17417 18748
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 2622 18652 2774 18680
rect 2746 18612 2774 18652
rect 5258 18640 5264 18692
rect 5316 18640 5322 18692
rect 5828 18652 6960 18680
rect 5828 18612 5856 18652
rect 2746 18584 5856 18612
rect 6932 18612 6960 18652
rect 7834 18640 7840 18692
rect 7892 18640 7898 18692
rect 8294 18680 8300 18692
rect 8255 18652 8300 18680
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 10410 18680 10416 18692
rect 8404 18652 10416 18680
rect 8404 18612 8432 18652
rect 10410 18640 10416 18652
rect 10468 18640 10474 18692
rect 11517 18683 11575 18689
rect 11517 18649 11529 18683
rect 11563 18649 11575 18683
rect 11517 18643 11575 18649
rect 12069 18683 12127 18689
rect 12069 18649 12081 18683
rect 12115 18680 12127 18683
rect 12158 18680 12164 18692
rect 12115 18652 12164 18680
rect 12115 18649 12127 18652
rect 12069 18643 12127 18649
rect 10134 18612 10140 18624
rect 6932 18584 8432 18612
rect 10095 18584 10140 18612
rect 10134 18572 10140 18584
rect 10192 18572 10198 18624
rect 10781 18615 10839 18621
rect 10781 18581 10793 18615
rect 10827 18612 10839 18615
rect 11532 18612 11560 18643
rect 12158 18640 12164 18652
rect 12216 18640 12222 18692
rect 12529 18683 12587 18689
rect 12529 18649 12541 18683
rect 12575 18649 12587 18683
rect 13078 18680 13084 18692
rect 13039 18652 13084 18680
rect 12529 18643 12587 18649
rect 10827 18584 11560 18612
rect 12544 18612 12572 18643
rect 13078 18640 13084 18652
rect 13136 18640 13142 18692
rect 13998 18640 14004 18692
rect 14056 18680 14062 18692
rect 14292 18680 14320 18708
rect 14829 18683 14887 18689
rect 14829 18680 14841 18683
rect 14056 18652 14841 18680
rect 14056 18640 14062 18652
rect 14829 18649 14841 18652
rect 14875 18649 14887 18683
rect 15378 18680 15384 18692
rect 15339 18652 15384 18680
rect 14829 18643 14887 18649
rect 15378 18640 15384 18652
rect 15436 18640 15442 18692
rect 17589 18683 17647 18689
rect 17589 18649 17601 18683
rect 17635 18680 17647 18683
rect 17954 18680 17960 18692
rect 17635 18652 17960 18680
rect 17635 18649 17647 18652
rect 17589 18643 17647 18649
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 18690 18680 18696 18692
rect 18651 18652 18696 18680
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 18782 18640 18788 18692
rect 18840 18680 18846 18692
rect 18840 18652 18885 18680
rect 18840 18640 18846 18652
rect 18966 18640 18972 18692
rect 19024 18680 19030 18692
rect 19613 18683 19671 18689
rect 19613 18680 19625 18683
rect 19024 18652 19625 18680
rect 19024 18640 19030 18652
rect 19613 18649 19625 18652
rect 19659 18649 19671 18683
rect 20533 18683 20591 18689
rect 20533 18680 20545 18683
rect 19613 18643 19671 18649
rect 19720 18652 20545 18680
rect 12618 18612 12624 18624
rect 12544 18584 12624 18612
rect 10827 18581 10839 18584
rect 10781 18575 10839 18581
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 15286 18572 15292 18624
rect 15344 18612 15350 18624
rect 19720 18612 19748 18652
rect 20533 18649 20545 18652
rect 20579 18680 20591 18683
rect 20622 18680 20628 18692
rect 20579 18652 20628 18680
rect 20579 18649 20591 18652
rect 20533 18643 20591 18649
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 21174 18680 21180 18692
rect 21135 18652 21180 18680
rect 21174 18640 21180 18652
rect 21232 18640 21238 18692
rect 21729 18683 21787 18689
rect 21729 18649 21741 18683
rect 21775 18649 21787 18683
rect 21729 18643 21787 18649
rect 15344 18584 19748 18612
rect 15344 18572 15350 18584
rect 19794 18572 19800 18624
rect 19852 18612 19858 18624
rect 21744 18612 21772 18643
rect 19852 18584 21772 18612
rect 19852 18572 19858 18584
rect 1104 18522 36892 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 36892 18522
rect 1104 18448 36892 18470
rect 1949 18411 2007 18417
rect 1949 18377 1961 18411
rect 1995 18408 2007 18411
rect 2498 18408 2504 18420
rect 1995 18380 2504 18408
rect 1995 18377 2007 18380
rect 1949 18371 2007 18377
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 5534 18408 5540 18420
rect 3476 18380 5540 18408
rect 3476 18368 3482 18380
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 6641 18411 6699 18417
rect 6641 18408 6653 18411
rect 6052 18380 6653 18408
rect 6052 18368 6058 18380
rect 6641 18377 6653 18380
rect 6687 18377 6699 18411
rect 10134 18408 10140 18420
rect 6641 18371 6699 18377
rect 7300 18380 10140 18408
rect 4338 18340 4344 18352
rect 2990 18312 4344 18340
rect 4338 18300 4344 18312
rect 4396 18300 4402 18352
rect 7300 18340 7328 18380
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 14366 18408 14372 18420
rect 10244 18380 14372 18408
rect 5198 18312 7328 18340
rect 7469 18343 7527 18349
rect 7469 18309 7481 18343
rect 7515 18340 7527 18343
rect 7558 18340 7564 18352
rect 7515 18312 7564 18340
rect 7515 18309 7527 18312
rect 7469 18303 7527 18309
rect 7558 18300 7564 18312
rect 7616 18300 7622 18352
rect 9766 18340 9772 18352
rect 8694 18312 9772 18340
rect 9766 18300 9772 18312
rect 9824 18300 9830 18352
rect 5902 18232 5908 18284
rect 5960 18272 5966 18284
rect 6733 18275 6791 18281
rect 5960 18244 6005 18272
rect 5960 18232 5966 18244
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 7006 18272 7012 18284
rect 6779 18244 7012 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 8846 18232 8852 18284
rect 8904 18272 8910 18284
rect 9858 18272 9864 18284
rect 8904 18244 9864 18272
rect 8904 18232 8910 18244
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 1946 18164 1952 18216
rect 2004 18164 2010 18216
rect 3418 18204 3424 18216
rect 3379 18176 3424 18204
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 3697 18207 3755 18213
rect 3697 18173 3709 18207
rect 3743 18204 3755 18207
rect 5626 18204 5632 18216
rect 3743 18176 4660 18204
rect 5587 18176 5632 18204
rect 3743 18173 3755 18176
rect 3697 18167 3755 18173
rect 1964 18136 1992 18164
rect 1964 18108 2452 18136
rect 2424 18068 2452 18108
rect 4157 18071 4215 18077
rect 4157 18068 4169 18071
rect 2424 18040 4169 18068
rect 4157 18037 4169 18040
rect 4203 18037 4215 18071
rect 4632 18068 4660 18176
rect 5626 18164 5632 18176
rect 5684 18164 5690 18216
rect 7190 18204 7196 18216
rect 5828 18176 7196 18204
rect 5828 18068 5856 18176
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 8754 18164 8760 18216
rect 8812 18204 8818 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 8812 18176 9229 18204
rect 8812 18164 8818 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 10244 18204 10272 18380
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 18693 18411 18751 18417
rect 18693 18377 18705 18411
rect 18739 18408 18751 18411
rect 18782 18408 18788 18420
rect 18739 18380 18788 18408
rect 18739 18377 18751 18380
rect 18693 18371 18751 18377
rect 18782 18368 18788 18380
rect 18840 18368 18846 18420
rect 21266 18408 21272 18420
rect 19352 18380 20668 18408
rect 21227 18380 21272 18408
rect 12066 18340 12072 18352
rect 12027 18312 12072 18340
rect 12066 18300 12072 18312
rect 12124 18300 12130 18352
rect 12618 18340 12624 18352
rect 12579 18312 12624 18340
rect 12618 18300 12624 18312
rect 12676 18300 12682 18352
rect 13722 18340 13728 18352
rect 13683 18312 13728 18340
rect 13722 18300 13728 18312
rect 13780 18300 13786 18352
rect 15194 18340 15200 18352
rect 15155 18312 15200 18340
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 15289 18343 15347 18349
rect 15289 18309 15301 18343
rect 15335 18340 15347 18343
rect 16945 18343 17003 18349
rect 16945 18340 16957 18343
rect 15335 18312 16957 18340
rect 15335 18309 15347 18312
rect 15289 18303 15347 18309
rect 16945 18309 16957 18312
rect 16991 18309 17003 18343
rect 16945 18303 17003 18309
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10410 18272 10416 18284
rect 10367 18244 10416 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 10870 18232 10876 18284
rect 10928 18272 10934 18284
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10928 18244 10977 18272
rect 10928 18232 10934 18244
rect 10965 18241 10977 18244
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 9364 18176 10272 18204
rect 11977 18207 12035 18213
rect 9364 18164 9370 18176
rect 11977 18173 11989 18207
rect 12023 18204 12035 18207
rect 12434 18204 12440 18216
rect 12023 18176 12440 18204
rect 12023 18173 12035 18176
rect 11977 18167 12035 18173
rect 12434 18164 12440 18176
rect 12492 18164 12498 18216
rect 8662 18096 8668 18148
rect 8720 18136 8726 18148
rect 12636 18136 12664 18300
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 16816 18244 17049 18272
rect 16816 18232 16822 18244
rect 17037 18241 17049 18244
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19352 18281 19380 18380
rect 19426 18300 19432 18352
rect 19484 18340 19490 18352
rect 20533 18343 20591 18349
rect 20533 18340 20545 18343
rect 19484 18312 20545 18340
rect 19484 18300 19490 18312
rect 20533 18309 20545 18312
rect 20579 18309 20591 18343
rect 20640 18340 20668 18380
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 22922 18408 22928 18420
rect 22883 18380 22928 18408
rect 22922 18368 22928 18380
rect 22980 18368 22986 18420
rect 27614 18340 27620 18352
rect 20640 18312 27620 18340
rect 20533 18303 20591 18309
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 19116 18244 19349 18272
rect 19116 18232 19122 18244
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 19337 18235 19395 18241
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 21361 18275 21419 18281
rect 21361 18272 21373 18275
rect 21140 18244 21373 18272
rect 21140 18232 21146 18244
rect 21361 18241 21373 18244
rect 21407 18241 21419 18275
rect 22462 18272 22468 18284
rect 22375 18244 22468 18272
rect 21361 18235 21419 18241
rect 22462 18232 22468 18244
rect 22520 18272 22526 18284
rect 22922 18272 22928 18284
rect 22520 18244 22928 18272
rect 22520 18232 22526 18244
rect 22922 18232 22928 18244
rect 22980 18232 22986 18284
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18272 25007 18275
rect 25501 18275 25559 18281
rect 25501 18272 25513 18275
rect 24995 18244 25513 18272
rect 24995 18241 25007 18244
rect 24949 18235 25007 18241
rect 25501 18241 25513 18244
rect 25547 18272 25559 18275
rect 34514 18272 34520 18284
rect 25547 18244 34520 18272
rect 25547 18241 25559 18244
rect 25501 18235 25559 18241
rect 34514 18232 34520 18244
rect 34572 18232 34578 18284
rect 36078 18272 36084 18284
rect 36039 18244 36084 18272
rect 36078 18232 36084 18244
rect 36136 18232 36142 18284
rect 13170 18164 13176 18216
rect 13228 18204 13234 18216
rect 13630 18204 13636 18216
rect 13228 18176 13636 18204
rect 13228 18164 13234 18176
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 14645 18207 14703 18213
rect 14645 18173 14657 18207
rect 14691 18204 14703 18207
rect 15286 18204 15292 18216
rect 14691 18176 15292 18204
rect 14691 18173 14703 18176
rect 14645 18167 14703 18173
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 15841 18207 15899 18213
rect 15841 18173 15853 18207
rect 15887 18204 15899 18207
rect 19242 18204 19248 18216
rect 15887 18176 19248 18204
rect 15887 18173 15899 18176
rect 15841 18167 15899 18173
rect 19242 18164 19248 18176
rect 19300 18164 19306 18216
rect 20162 18204 20168 18216
rect 20123 18176 20168 18204
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 20622 18204 20628 18216
rect 20583 18176 20628 18204
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 8720 18108 12664 18136
rect 8720 18096 8726 18108
rect 21726 18096 21732 18148
rect 21784 18136 21790 18148
rect 24857 18139 24915 18145
rect 24857 18136 24869 18139
rect 21784 18108 24869 18136
rect 21784 18096 21790 18108
rect 24857 18105 24869 18108
rect 24903 18105 24915 18139
rect 24857 18099 24915 18105
rect 4632 18040 5856 18068
rect 4157 18031 4215 18037
rect 6178 18028 6184 18080
rect 6236 18068 6242 18080
rect 10229 18071 10287 18077
rect 10229 18068 10241 18071
rect 6236 18040 10241 18068
rect 6236 18028 6242 18040
rect 10229 18037 10241 18040
rect 10275 18037 10287 18071
rect 10229 18031 10287 18037
rect 11057 18071 11115 18077
rect 11057 18037 11069 18071
rect 11103 18068 11115 18071
rect 11974 18068 11980 18080
rect 11103 18040 11980 18068
rect 11103 18037 11115 18040
rect 11057 18031 11115 18037
rect 11974 18028 11980 18040
rect 12032 18028 12038 18080
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 17954 18068 17960 18080
rect 17911 18040 17960 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 17954 18028 17960 18040
rect 18012 18068 18018 18080
rect 19334 18068 19340 18080
rect 18012 18040 19340 18068
rect 18012 18028 18018 18040
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 19429 18071 19487 18077
rect 19429 18037 19441 18071
rect 19475 18068 19487 18071
rect 19978 18068 19984 18080
rect 19475 18040 19984 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 22370 18068 22376 18080
rect 22331 18040 22376 18068
rect 22370 18028 22376 18040
rect 22428 18028 22434 18080
rect 36262 18068 36268 18080
rect 36223 18040 36268 18068
rect 36262 18028 36268 18040
rect 36320 18028 36326 18080
rect 1104 17978 36892 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 36892 17978
rect 1104 17904 36892 17926
rect 1844 17867 1902 17873
rect 1844 17833 1856 17867
rect 1890 17864 1902 17867
rect 8478 17864 8484 17876
rect 1890 17836 4476 17864
rect 8439 17836 8484 17864
rect 1890 17833 1902 17836
rect 1844 17827 1902 17833
rect 3329 17799 3387 17805
rect 3329 17765 3341 17799
rect 3375 17796 3387 17799
rect 3510 17796 3516 17808
rect 3375 17768 3516 17796
rect 3375 17765 3387 17768
rect 3329 17759 3387 17765
rect 3510 17756 3516 17768
rect 3568 17756 3574 17808
rect 4448 17796 4476 17836
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 10778 17864 10784 17876
rect 10739 17836 10784 17864
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 12526 17824 12532 17876
rect 12584 17864 12590 17876
rect 16117 17867 16175 17873
rect 12584 17836 16068 17864
rect 12584 17824 12590 17836
rect 4448 17768 4568 17796
rect 2406 17688 2412 17740
rect 2464 17728 2470 17740
rect 4062 17728 4068 17740
rect 2464 17700 4068 17728
rect 2464 17688 2470 17700
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 4430 17728 4436 17740
rect 4391 17700 4436 17728
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 4540 17728 4568 17768
rect 6730 17756 6736 17808
rect 6788 17756 6794 17808
rect 8110 17756 8116 17808
rect 8168 17796 8174 17808
rect 9493 17799 9551 17805
rect 9493 17796 9505 17799
rect 8168 17768 9505 17796
rect 8168 17756 8174 17768
rect 9493 17765 9505 17768
rect 9539 17765 9551 17799
rect 9493 17759 9551 17765
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 16040 17796 16068 17836
rect 16117 17833 16129 17867
rect 16163 17864 16175 17867
rect 19426 17864 19432 17876
rect 16163 17836 19432 17864
rect 16163 17833 16175 17836
rect 16117 17827 16175 17833
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 21913 17867 21971 17873
rect 21913 17833 21925 17867
rect 21959 17864 21971 17867
rect 22094 17864 22100 17876
rect 21959 17836 22100 17864
rect 21959 17833 21971 17836
rect 21913 17827 21971 17833
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 10928 17768 15332 17796
rect 16040 17768 16160 17796
rect 10928 17756 10934 17768
rect 6362 17728 6368 17740
rect 4540 17700 6368 17728
rect 6362 17688 6368 17700
rect 6420 17688 6426 17740
rect 6454 17688 6460 17740
rect 6512 17728 6518 17740
rect 6748 17728 6776 17756
rect 7009 17731 7067 17737
rect 7009 17728 7021 17731
rect 6512 17700 7021 17728
rect 6512 17688 6518 17700
rect 7009 17697 7021 17700
rect 7055 17697 7067 17731
rect 7009 17691 7067 17697
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 10137 17731 10195 17737
rect 10137 17728 10149 17731
rect 7800 17700 10149 17728
rect 7800 17688 7806 17700
rect 10137 17697 10149 17700
rect 10183 17697 10195 17731
rect 10137 17691 10195 17697
rect 10502 17688 10508 17740
rect 10560 17728 10566 17740
rect 11517 17731 11575 17737
rect 11517 17728 11529 17731
rect 10560 17700 11529 17728
rect 10560 17688 10566 17700
rect 11517 17697 11529 17700
rect 11563 17697 11575 17731
rect 11517 17691 11575 17697
rect 12158 17688 12164 17740
rect 12216 17728 12222 17740
rect 12216 17700 12434 17728
rect 12216 17688 12222 17700
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 6733 17663 6791 17669
rect 6733 17629 6745 17663
rect 6779 17629 6791 17663
rect 6733 17623 6791 17629
rect 3082 17564 4660 17592
rect 4632 17524 4660 17564
rect 4706 17552 4712 17604
rect 4764 17592 4770 17604
rect 6638 17592 6644 17604
rect 4764 17564 5120 17592
rect 5934 17564 6644 17592
rect 4764 17552 4770 17564
rect 4798 17524 4804 17536
rect 4632 17496 4804 17524
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 5092 17524 5120 17564
rect 6638 17552 6644 17564
rect 6696 17552 6702 17604
rect 6748 17592 6776 17623
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9582 17660 9588 17672
rect 8904 17632 9588 17660
rect 8904 17620 8910 17632
rect 9582 17620 9588 17632
rect 9640 17660 9646 17672
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 9640 17632 10241 17660
rect 9640 17620 9646 17632
rect 10229 17629 10241 17632
rect 10275 17660 10287 17663
rect 10410 17660 10416 17672
rect 10275 17632 10416 17660
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 10594 17620 10600 17672
rect 10652 17660 10658 17672
rect 10873 17663 10931 17669
rect 10873 17660 10885 17663
rect 10652 17632 10885 17660
rect 10652 17620 10658 17632
rect 10873 17629 10885 17632
rect 10919 17629 10931 17663
rect 12406 17660 12434 17700
rect 13262 17688 13268 17740
rect 13320 17728 13326 17740
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 13320 17700 13369 17728
rect 13320 17688 13326 17700
rect 13357 17697 13369 17700
rect 13403 17728 13415 17731
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13403 17700 14289 17728
rect 13403 17697 13415 17700
rect 13357 17691 13415 17697
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 14921 17731 14979 17737
rect 14921 17697 14933 17731
rect 14967 17728 14979 17731
rect 15194 17728 15200 17740
rect 14967 17700 15200 17728
rect 14967 17697 14979 17700
rect 14921 17691 14979 17697
rect 15194 17688 15200 17700
rect 15252 17688 15258 17740
rect 15304 17728 15332 17768
rect 15304 17700 16068 17728
rect 12710 17660 12716 17672
rect 12406 17632 12716 17660
rect 10873 17623 10931 17629
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 16040 17669 16068 17700
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17629 16083 17663
rect 16132 17660 16160 17768
rect 16758 17756 16764 17808
rect 16816 17796 16822 17808
rect 17313 17799 17371 17805
rect 17313 17796 17325 17799
rect 16816 17768 17325 17796
rect 16816 17756 16822 17768
rect 17313 17765 17325 17768
rect 17359 17765 17371 17799
rect 17313 17759 17371 17765
rect 20162 17756 20168 17808
rect 20220 17796 20226 17808
rect 22370 17796 22376 17808
rect 20220 17768 21220 17796
rect 20220 17756 20226 17768
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 20530 17728 20536 17740
rect 16448 17700 18184 17728
rect 20491 17700 20536 17728
rect 16448 17688 16454 17700
rect 16669 17663 16727 17669
rect 16669 17660 16681 17663
rect 16132 17632 16681 17660
rect 16025 17623 16083 17629
rect 16669 17629 16681 17632
rect 16715 17629 16727 17663
rect 16669 17623 16727 17629
rect 7282 17592 7288 17604
rect 6748 17564 7288 17592
rect 7282 17552 7288 17564
rect 7340 17552 7346 17604
rect 9674 17592 9680 17604
rect 8234 17564 9680 17592
rect 9674 17552 9680 17564
rect 9732 17552 9738 17604
rect 11606 17552 11612 17604
rect 11664 17592 11670 17604
rect 12161 17595 12219 17601
rect 11664 17564 11709 17592
rect 11664 17552 11670 17564
rect 12161 17561 12173 17595
rect 12207 17592 12219 17595
rect 12618 17592 12624 17604
rect 12207 17564 12624 17592
rect 12207 17561 12219 17564
rect 12161 17555 12219 17561
rect 12618 17552 12624 17564
rect 12676 17552 12682 17604
rect 13078 17592 13084 17604
rect 13039 17564 13084 17592
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 13173 17595 13231 17601
rect 13173 17561 13185 17595
rect 13219 17561 13231 17595
rect 14826 17592 14832 17604
rect 14787 17564 14832 17592
rect 13173 17555 13231 17561
rect 5718 17524 5724 17536
rect 5092 17496 5724 17524
rect 5718 17484 5724 17496
rect 5776 17484 5782 17536
rect 6181 17527 6239 17533
rect 6181 17493 6193 17527
rect 6227 17524 6239 17527
rect 7650 17524 7656 17536
rect 6227 17496 7656 17524
rect 6227 17493 6239 17496
rect 6181 17487 6239 17493
rect 7650 17484 7656 17496
rect 7708 17524 7714 17536
rect 10042 17524 10048 17536
rect 7708 17496 10048 17524
rect 7708 17484 7714 17496
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 12434 17484 12440 17536
rect 12492 17524 12498 17536
rect 13096 17524 13124 17552
rect 12492 17496 13124 17524
rect 13188 17524 13216 17555
rect 14826 17552 14832 17564
rect 14884 17552 14890 17604
rect 18156 17601 18184 17700
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 21192 17737 21220 17768
rect 21560 17768 22376 17796
rect 21177 17731 21235 17737
rect 21177 17697 21189 17731
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 19426 17620 19432 17672
rect 19484 17660 19490 17672
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 19484 17632 19625 17660
rect 19484 17620 19490 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 16761 17595 16819 17601
rect 16761 17592 16773 17595
rect 15028 17564 16773 17592
rect 15028 17524 15056 17564
rect 16761 17561 16773 17564
rect 16807 17561 16819 17595
rect 16761 17555 16819 17561
rect 18141 17595 18199 17601
rect 18141 17561 18153 17595
rect 18187 17592 18199 17595
rect 18230 17592 18236 17604
rect 18187 17564 18236 17592
rect 18187 17561 18199 17564
rect 18141 17555 18199 17561
rect 18230 17552 18236 17564
rect 18288 17592 18294 17604
rect 20990 17592 20996 17604
rect 18288 17564 20996 17592
rect 18288 17552 18294 17564
rect 20990 17552 20996 17564
rect 21048 17552 21054 17604
rect 21085 17595 21143 17601
rect 21085 17561 21097 17595
rect 21131 17561 21143 17595
rect 21085 17555 21143 17561
rect 13188 17496 15056 17524
rect 15565 17527 15623 17533
rect 12492 17484 12498 17496
rect 15565 17493 15577 17527
rect 15611 17524 15623 17527
rect 15930 17524 15936 17536
rect 15611 17496 15936 17524
rect 15611 17493 15623 17496
rect 15565 17487 15623 17493
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 18877 17527 18935 17533
rect 18877 17493 18889 17527
rect 18923 17524 18935 17527
rect 19058 17524 19064 17536
rect 18923 17496 19064 17524
rect 18923 17493 18935 17496
rect 18877 17487 18935 17493
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 19521 17527 19579 17533
rect 19521 17493 19533 17527
rect 19567 17524 19579 17527
rect 20162 17524 20168 17536
rect 19567 17496 20168 17524
rect 19567 17493 19579 17496
rect 19521 17487 19579 17493
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 21100 17524 21128 17555
rect 21560 17524 21588 17768
rect 22370 17756 22376 17768
rect 22428 17756 22434 17808
rect 21634 17688 21640 17740
rect 21692 17728 21698 17740
rect 23017 17731 23075 17737
rect 23017 17728 23029 17731
rect 21692 17700 23029 17728
rect 21692 17688 21698 17700
rect 23017 17697 23029 17700
rect 23063 17697 23075 17731
rect 23017 17691 23075 17697
rect 21818 17660 21824 17672
rect 21731 17632 21824 17660
rect 21818 17620 21824 17632
rect 21876 17660 21882 17672
rect 21876 17632 22600 17660
rect 21876 17620 21882 17632
rect 22572 17601 22600 17632
rect 22557 17595 22615 17601
rect 22557 17561 22569 17595
rect 22603 17592 22615 17595
rect 22603 17564 26234 17592
rect 22603 17561 22615 17564
rect 22557 17555 22615 17561
rect 21100 17496 21588 17524
rect 26206 17524 26234 17564
rect 36538 17524 36544 17536
rect 26206 17496 36544 17524
rect 36538 17484 36544 17496
rect 36596 17484 36602 17536
rect 1104 17434 36892 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 36892 17434
rect 1104 17360 36892 17382
rect 1670 17320 1676 17332
rect 1631 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 3970 17280 3976 17332
rect 4028 17320 4034 17332
rect 4801 17323 4859 17329
rect 4028 17292 4660 17320
rect 4028 17280 4034 17292
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 1636 17224 2774 17252
rect 1636 17212 1642 17224
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 1857 17187 1915 17193
rect 1857 17184 1869 17187
rect 1544 17156 1869 17184
rect 1544 17144 1550 17156
rect 1857 17153 1869 17156
rect 1903 17153 1915 17187
rect 1857 17147 1915 17153
rect 2593 17187 2651 17193
rect 2593 17153 2605 17187
rect 2639 17153 2651 17187
rect 2593 17147 2651 17153
rect 2406 17048 2412 17060
rect 2367 17020 2412 17048
rect 2406 17008 2412 17020
rect 2464 17008 2470 17060
rect 2608 17048 2636 17147
rect 2746 17116 2774 17224
rect 3786 17212 3792 17264
rect 3844 17212 3850 17264
rect 4632 17252 4660 17292
rect 4801 17289 4813 17323
rect 4847 17320 4859 17323
rect 5534 17320 5540 17332
rect 4847 17292 5540 17320
rect 4847 17289 4859 17292
rect 4801 17283 4859 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 6638 17280 6644 17332
rect 6696 17320 6702 17332
rect 6733 17323 6791 17329
rect 6733 17320 6745 17323
rect 6696 17292 6745 17320
rect 6696 17280 6702 17292
rect 6733 17289 6745 17292
rect 6779 17289 6791 17323
rect 6733 17283 6791 17289
rect 6840 17292 9674 17320
rect 6840 17252 6868 17292
rect 4632 17224 6868 17252
rect 7098 17212 7104 17264
rect 7156 17252 7162 17264
rect 7561 17255 7619 17261
rect 7561 17252 7573 17255
rect 7156 17224 7573 17252
rect 7156 17212 7162 17224
rect 7561 17221 7573 17224
rect 7607 17252 7619 17255
rect 7834 17252 7840 17264
rect 7607 17224 7840 17252
rect 7607 17221 7619 17224
rect 7561 17215 7619 17221
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 9214 17252 9220 17264
rect 8786 17224 9220 17252
rect 9214 17212 9220 17224
rect 9272 17212 9278 17264
rect 5994 17184 6000 17196
rect 5955 17156 6000 17184
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 6270 17144 6276 17196
rect 6328 17184 6334 17196
rect 6822 17184 6828 17196
rect 6328 17156 6828 17184
rect 6328 17144 6334 17156
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 3053 17119 3111 17125
rect 3053 17116 3065 17119
rect 2746 17088 3065 17116
rect 3053 17085 3065 17088
rect 3099 17116 3111 17119
rect 3329 17119 3387 17125
rect 3099 17088 3188 17116
rect 3099 17085 3111 17088
rect 3053 17079 3111 17085
rect 2958 17048 2964 17060
rect 2608 17020 2964 17048
rect 2958 17008 2964 17020
rect 3016 17008 3022 17060
rect 3160 16980 3188 17088
rect 3329 17085 3341 17119
rect 3375 17116 3387 17119
rect 3694 17116 3700 17128
rect 3375 17088 3700 17116
rect 3375 17085 3387 17088
rect 3329 17079 3387 17085
rect 3694 17076 3700 17088
rect 3752 17076 3758 17128
rect 3970 17076 3976 17128
rect 4028 17116 4034 17128
rect 7282 17116 7288 17128
rect 4028 17088 7144 17116
rect 7243 17088 7288 17116
rect 4028 17076 4034 17088
rect 7116 17048 7144 17088
rect 7282 17076 7288 17088
rect 7340 17076 7346 17128
rect 9309 17119 9367 17125
rect 9309 17116 9321 17119
rect 7392 17088 9321 17116
rect 7392 17048 7420 17088
rect 9309 17085 9321 17088
rect 9355 17085 9367 17119
rect 9646 17116 9674 17292
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10321 17323 10379 17329
rect 10321 17320 10333 17323
rect 10284 17292 10333 17320
rect 10284 17280 10290 17292
rect 10321 17289 10333 17292
rect 10367 17289 10379 17323
rect 10321 17283 10379 17289
rect 10410 17280 10416 17332
rect 10468 17280 10474 17332
rect 11057 17323 11115 17329
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 11606 17320 11612 17332
rect 11103 17292 11612 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 21634 17320 21640 17332
rect 11707 17292 21640 17320
rect 10428 17252 10456 17280
rect 11707 17252 11735 17292
rect 21634 17280 21640 17292
rect 21692 17280 21698 17332
rect 11882 17252 11888 17264
rect 10428 17224 11735 17252
rect 11843 17224 11888 17252
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 11974 17212 11980 17264
rect 12032 17252 12038 17264
rect 13081 17255 13139 17261
rect 13081 17252 13093 17255
rect 12032 17224 13093 17252
rect 12032 17212 12038 17224
rect 13081 17221 13093 17224
rect 13127 17221 13139 17255
rect 13081 17215 13139 17221
rect 13630 17212 13636 17264
rect 13688 17252 13694 17264
rect 14829 17255 14887 17261
rect 14829 17252 14841 17255
rect 13688 17224 14841 17252
rect 13688 17212 13694 17224
rect 14829 17221 14841 17224
rect 14875 17221 14887 17255
rect 14829 17215 14887 17221
rect 15378 17212 15384 17264
rect 15436 17252 15442 17264
rect 16390 17252 16396 17264
rect 15436 17224 15481 17252
rect 16132 17224 16396 17252
rect 15436 17212 15442 17224
rect 10410 17184 10416 17196
rect 10371 17156 10416 17184
rect 10410 17144 10416 17156
rect 10468 17144 10474 17196
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17184 11023 17187
rect 11146 17184 11152 17196
rect 11011 17156 11152 17184
rect 11011 17153 11023 17156
rect 10965 17147 11023 17153
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17184 14427 17187
rect 16132 17184 16160 17224
rect 16390 17212 16396 17224
rect 16448 17212 16454 17264
rect 17494 17212 17500 17264
rect 17552 17252 17558 17264
rect 20441 17255 20499 17261
rect 20441 17252 20453 17255
rect 17552 17224 20453 17252
rect 17552 17212 17558 17224
rect 20441 17221 20453 17224
rect 20487 17221 20499 17255
rect 20990 17252 20996 17264
rect 20951 17224 20996 17252
rect 20441 17215 20499 17221
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 21082 17212 21088 17264
rect 21140 17252 21146 17264
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21140 17224 22017 17252
rect 21140 17212 21146 17224
rect 22005 17221 22017 17224
rect 22051 17221 22063 17255
rect 22005 17215 22063 17221
rect 14415 17156 14872 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 11793 17119 11851 17125
rect 9646 17088 11744 17116
rect 9309 17079 9367 17085
rect 7116 17020 7420 17048
rect 9324 17048 9352 17079
rect 11716 17048 11744 17088
rect 11793 17085 11805 17119
rect 11839 17116 11851 17119
rect 12158 17116 12164 17128
rect 11839 17088 12164 17116
rect 11839 17085 11851 17088
rect 11793 17079 11851 17085
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 12986 17116 12992 17128
rect 12268 17088 12992 17116
rect 12268 17048 12296 17088
rect 12986 17076 12992 17088
rect 13044 17076 13050 17128
rect 13633 17119 13691 17125
rect 13633 17085 13645 17119
rect 13679 17116 13691 17119
rect 14090 17116 14096 17128
rect 13679 17088 14096 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 9324 17020 10824 17048
rect 11716 17020 12296 17048
rect 12345 17051 12403 17057
rect 4430 16980 4436 16992
rect 3160 16952 4436 16980
rect 4430 16940 4436 16952
rect 4488 16980 4494 16992
rect 4706 16980 4712 16992
rect 4488 16952 4712 16980
rect 4488 16940 4494 16952
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 5905 16983 5963 16989
rect 5905 16980 5917 16983
rect 5592 16952 5917 16980
rect 5592 16940 5598 16952
rect 5905 16949 5917 16952
rect 5951 16949 5963 16983
rect 5905 16943 5963 16949
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 10686 16980 10692 16992
rect 7432 16952 10692 16980
rect 7432 16940 7438 16952
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 10796 16980 10824 17020
rect 12345 17017 12357 17051
rect 12391 17048 12403 17051
rect 13262 17048 13268 17060
rect 12391 17020 13268 17048
rect 12391 17017 12403 17020
rect 12345 17011 12403 17017
rect 13262 17008 13268 17020
rect 13320 17008 13326 17060
rect 14384 17048 14412 17147
rect 14108 17020 14412 17048
rect 14844 17048 14872 17156
rect 15672 17156 16160 17184
rect 16209 17187 16267 17193
rect 15102 17076 15108 17128
rect 15160 17116 15166 17128
rect 15473 17119 15531 17125
rect 15473 17116 15485 17119
rect 15160 17088 15485 17116
rect 15160 17076 15166 17088
rect 15473 17085 15485 17088
rect 15519 17085 15531 17119
rect 15473 17079 15531 17085
rect 15672 17048 15700 17156
rect 16209 17153 16221 17187
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 17773 17187 17831 17193
rect 17773 17153 17785 17187
rect 17819 17184 17831 17187
rect 18417 17187 18475 17193
rect 18417 17184 18429 17187
rect 17819 17156 18429 17184
rect 17819 17153 17831 17156
rect 17773 17147 17831 17153
rect 18417 17153 18429 17156
rect 18463 17184 18475 17187
rect 19061 17187 19119 17193
rect 19061 17184 19073 17187
rect 18463 17156 19073 17184
rect 18463 17153 18475 17156
rect 18417 17147 18475 17153
rect 19061 17153 19073 17156
rect 19107 17184 19119 17187
rect 19107 17156 19840 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 16224 17116 16252 17147
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 14844 17020 15700 17048
rect 15764 17088 16865 17116
rect 14108 16980 14136 17020
rect 14274 16980 14280 16992
rect 10796 16952 14136 16980
rect 14235 16952 14280 16980
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15764 16980 15792 17088
rect 16853 17085 16865 17088
rect 16899 17116 16911 17119
rect 19610 17116 19616 17128
rect 16899 17088 19616 17116
rect 16899 17085 16911 17088
rect 16853 17079 16911 17085
rect 19610 17076 19616 17088
rect 19668 17076 19674 17128
rect 16390 17008 16396 17060
rect 16448 17048 16454 17060
rect 18414 17048 18420 17060
rect 16448 17020 18420 17048
rect 16448 17008 16454 17020
rect 18414 17008 18420 17020
rect 18472 17008 18478 17060
rect 18874 17048 18880 17060
rect 18835 17020 18880 17048
rect 18874 17008 18880 17020
rect 18932 17008 18938 17060
rect 19812 16992 19840 17156
rect 21085 17119 21143 17125
rect 21085 17085 21097 17119
rect 21131 17116 21143 17119
rect 21726 17116 21732 17128
rect 21131 17088 21732 17116
rect 21131 17085 21143 17088
rect 21085 17079 21143 17085
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 21450 17008 21456 17060
rect 21508 17048 21514 17060
rect 21508 17020 22094 17048
rect 21508 17008 21514 17020
rect 15068 16952 15792 16980
rect 15068 16940 15074 16952
rect 15838 16940 15844 16992
rect 15896 16980 15902 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 15896 16952 16129 16980
rect 15896 16940 15902 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 18322 16980 18328 16992
rect 18283 16952 18328 16980
rect 16117 16943 16175 16949
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19702 16980 19708 16992
rect 19484 16952 19708 16980
rect 19484 16940 19490 16952
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 19794 16940 19800 16992
rect 19852 16980 19858 16992
rect 21542 16980 21548 16992
rect 19852 16952 21548 16980
rect 19852 16940 19858 16952
rect 21542 16940 21548 16952
rect 21600 16940 21606 16992
rect 22066 16980 22094 17020
rect 22462 16980 22468 16992
rect 22066 16952 22468 16980
rect 22462 16940 22468 16952
rect 22520 16940 22526 16992
rect 1104 16890 36892 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 36892 16890
rect 1104 16816 36892 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1854 16776 1860 16788
rect 1728 16748 1860 16776
rect 1728 16736 1734 16748
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 3326 16776 3332 16788
rect 3287 16748 3332 16776
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 4120 16748 12434 16776
rect 4120 16736 4126 16748
rect 7285 16711 7343 16717
rect 7285 16677 7297 16711
rect 7331 16708 7343 16711
rect 7374 16708 7380 16720
rect 7331 16680 7380 16708
rect 7331 16677 7343 16680
rect 7285 16671 7343 16677
rect 7374 16668 7380 16680
rect 7432 16668 7438 16720
rect 7742 16668 7748 16720
rect 7800 16708 7806 16720
rect 12406 16708 12434 16748
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 18966 16776 18972 16788
rect 12584 16748 18972 16776
rect 12584 16736 12590 16748
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19521 16779 19579 16785
rect 19521 16745 19533 16779
rect 19567 16776 19579 16779
rect 19794 16776 19800 16788
rect 19567 16748 19800 16776
rect 19567 16745 19579 16748
rect 19521 16739 19579 16745
rect 19794 16736 19800 16748
rect 19852 16736 19858 16788
rect 20809 16779 20867 16785
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 20990 16776 20996 16788
rect 20855 16748 20996 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 21450 16776 21456 16788
rect 21411 16748 21456 16776
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 21542 16736 21548 16788
rect 21600 16776 21606 16788
rect 21600 16748 26234 16776
rect 21600 16736 21606 16748
rect 17405 16711 17463 16717
rect 7800 16680 11376 16708
rect 12406 16680 13216 16708
rect 7800 16668 7806 16680
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 3142 16600 3148 16652
rect 3200 16640 3206 16652
rect 3970 16640 3976 16652
rect 3200 16612 3976 16640
rect 3200 16600 3206 16612
rect 3970 16600 3976 16612
rect 4028 16600 4034 16652
rect 4246 16640 4252 16652
rect 4207 16612 4252 16640
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 4706 16640 4712 16652
rect 4619 16612 4712 16640
rect 4706 16600 4712 16612
rect 4764 16640 4770 16652
rect 9125 16643 9183 16649
rect 9125 16640 9137 16643
rect 4764 16612 9137 16640
rect 4764 16600 4770 16612
rect 9125 16609 9137 16612
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 6730 16572 6736 16584
rect 6691 16544 6736 16572
rect 6730 16532 6736 16544
rect 6788 16532 6794 16584
rect 7006 16532 7012 16584
rect 7064 16572 7070 16584
rect 7926 16572 7932 16584
rect 7064 16544 7932 16572
rect 7064 16532 7070 16544
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 8202 16532 8208 16584
rect 8260 16572 8266 16584
rect 8481 16575 8539 16581
rect 8481 16572 8493 16575
rect 8260 16544 8493 16572
rect 8260 16532 8266 16544
rect 8481 16541 8493 16544
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 8846 16572 8852 16584
rect 8619 16544 8852 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8846 16532 8852 16544
rect 8904 16532 8910 16584
rect 11348 16581 11376 16680
rect 13188 16652 13216 16680
rect 17405 16677 17417 16711
rect 17451 16708 17463 16711
rect 18046 16708 18052 16720
rect 17451 16680 18052 16708
rect 17451 16677 17463 16680
rect 17405 16671 17463 16677
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 19702 16668 19708 16720
rect 19760 16708 19766 16720
rect 20346 16708 20352 16720
rect 19760 16680 20352 16708
rect 19760 16668 19766 16680
rect 20346 16668 20352 16680
rect 20404 16668 20410 16720
rect 21468 16708 21496 16736
rect 21910 16708 21916 16720
rect 20732 16680 21496 16708
rect 21871 16680 21916 16708
rect 11425 16643 11483 16649
rect 11425 16609 11437 16643
rect 11471 16640 11483 16643
rect 12526 16640 12532 16652
rect 11471 16612 12532 16640
rect 11471 16609 11483 16612
rect 11425 16603 11483 16609
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 13170 16640 13176 16652
rect 13131 16612 13176 16640
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 15654 16640 15660 16652
rect 15615 16612 15660 16640
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 15979 16612 16865 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16853 16609 16865 16612
rect 16899 16640 16911 16643
rect 18322 16640 18328 16652
rect 16899 16612 18328 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 18322 16600 18328 16612
rect 18380 16600 18386 16652
rect 19610 16600 19616 16652
rect 19668 16640 19674 16652
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19668 16612 19993 16640
rect 19668 16600 19674 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12207 16544 12434 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 4890 16504 4896 16516
rect 3082 16476 4896 16504
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 4985 16507 5043 16513
rect 4985 16473 4997 16507
rect 5031 16504 5043 16507
rect 5074 16504 5080 16516
rect 5031 16476 5080 16504
rect 5031 16473 5043 16476
rect 4985 16467 5043 16473
rect 5074 16464 5080 16476
rect 5132 16464 5138 16516
rect 5718 16464 5724 16516
rect 5776 16464 5782 16516
rect 10873 16507 10931 16513
rect 10873 16504 10885 16507
rect 6656 16476 10885 16504
rect 4522 16396 4528 16448
rect 4580 16436 4586 16448
rect 5166 16436 5172 16448
rect 4580 16408 5172 16436
rect 4580 16396 4586 16408
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 5350 16396 5356 16448
rect 5408 16436 5414 16448
rect 6656 16436 6684 16476
rect 10873 16473 10885 16476
rect 10919 16504 10931 16507
rect 12406 16504 12434 16544
rect 14642 16532 14648 16584
rect 14700 16572 14706 16584
rect 14829 16575 14887 16581
rect 14829 16572 14841 16575
rect 14700 16544 14841 16572
rect 14700 16532 14706 16544
rect 14829 16541 14841 16544
rect 14875 16541 14887 16575
rect 18230 16572 18236 16584
rect 18191 16544 18236 16572
rect 14829 16535 14887 16541
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 20530 16572 20536 16584
rect 18564 16544 20536 16572
rect 18564 16532 18570 16544
rect 20530 16532 20536 16544
rect 20588 16532 20594 16584
rect 20732 16581 20760 16680
rect 21910 16668 21916 16680
rect 21968 16668 21974 16720
rect 22465 16711 22523 16717
rect 22465 16708 22477 16711
rect 22066 16680 22477 16708
rect 22066 16640 22094 16680
rect 22465 16677 22477 16680
rect 22511 16677 22523 16711
rect 26206 16708 26234 16748
rect 36446 16708 36452 16720
rect 26206 16680 36452 16708
rect 22465 16671 22523 16677
rect 36446 16668 36452 16680
rect 36504 16668 36510 16720
rect 20824 16612 22094 16640
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 12713 16507 12771 16513
rect 12713 16504 12725 16507
rect 10919 16476 11560 16504
rect 12406 16476 12725 16504
rect 10919 16473 10931 16476
rect 10873 16467 10931 16473
rect 5408 16408 6684 16436
rect 5408 16396 5414 16408
rect 7374 16396 7380 16448
rect 7432 16436 7438 16448
rect 7837 16439 7895 16445
rect 7837 16436 7849 16439
rect 7432 16408 7849 16436
rect 7432 16396 7438 16408
rect 7837 16405 7849 16408
rect 7883 16405 7895 16439
rect 7837 16399 7895 16405
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 11238 16436 11244 16448
rect 10836 16408 11244 16436
rect 10836 16396 10842 16408
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 11532 16436 11560 16476
rect 12713 16473 12725 16476
rect 12759 16473 12771 16507
rect 12713 16467 12771 16473
rect 12805 16507 12863 16513
rect 12805 16473 12817 16507
rect 12851 16504 12863 16507
rect 14274 16504 14280 16516
rect 12851 16476 14280 16504
rect 12851 16473 12863 16476
rect 12805 16467 12863 16473
rect 14274 16464 14280 16476
rect 14332 16464 14338 16516
rect 15838 16504 15844 16516
rect 14568 16476 14872 16504
rect 15799 16476 15844 16504
rect 14568 16436 14596 16476
rect 11532 16408 14596 16436
rect 14642 16396 14648 16448
rect 14700 16436 14706 16448
rect 14844 16436 14872 16476
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 20824 16504 20852 16612
rect 17000 16476 17045 16504
rect 17236 16476 20852 16504
rect 17000 16464 17006 16476
rect 17236 16436 17264 16476
rect 14700 16408 14745 16436
rect 14844 16408 17264 16436
rect 18325 16439 18383 16445
rect 14700 16396 14706 16408
rect 18325 16405 18337 16439
rect 18371 16436 18383 16439
rect 19334 16436 19340 16448
rect 18371 16408 19340 16436
rect 18371 16405 18383 16408
rect 18325 16399 18383 16405
rect 19334 16396 19340 16408
rect 19392 16396 19398 16448
rect 1104 16346 36892 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 36892 16346
rect 1104 16272 36892 16294
rect 4890 16192 4896 16244
rect 4948 16232 4954 16244
rect 6914 16232 6920 16244
rect 4948 16204 6920 16232
rect 4948 16192 4954 16204
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 9030 16232 9036 16244
rect 7300 16204 9036 16232
rect 2869 16167 2927 16173
rect 2869 16133 2881 16167
rect 2915 16164 2927 16167
rect 3234 16164 3240 16176
rect 2915 16136 3240 16164
rect 2915 16133 2927 16136
rect 2869 16127 2927 16133
rect 3234 16124 3240 16136
rect 3292 16124 3298 16176
rect 4186 16136 5304 16164
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 2682 16096 2688 16108
rect 1903 16068 2688 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 4893 16099 4951 16105
rect 4893 16065 4905 16099
rect 4939 16096 4951 16099
rect 4982 16096 4988 16108
rect 4939 16068 4988 16096
rect 4939 16065 4951 16068
rect 4893 16059 4951 16065
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 5276 16096 5304 16136
rect 6730 16124 6736 16176
rect 6788 16164 6794 16176
rect 7300 16164 7328 16204
rect 9030 16192 9036 16204
rect 9088 16232 9094 16244
rect 11885 16235 11943 16241
rect 9088 16204 11836 16232
rect 9088 16192 9094 16204
rect 6788 16136 7328 16164
rect 6788 16124 6794 16136
rect 7374 16124 7380 16176
rect 7432 16124 7438 16176
rect 7650 16164 7656 16176
rect 7611 16136 7656 16164
rect 7650 16124 7656 16136
rect 7708 16124 7714 16176
rect 9306 16164 9312 16176
rect 8878 16136 9312 16164
rect 9306 16124 9312 16136
rect 9364 16124 9370 16176
rect 10137 16167 10195 16173
rect 10137 16133 10149 16167
rect 10183 16164 10195 16167
rect 10226 16164 10232 16176
rect 10183 16136 10232 16164
rect 10183 16133 10195 16136
rect 10137 16127 10195 16133
rect 10226 16124 10232 16136
rect 10284 16164 10290 16176
rect 10686 16164 10692 16176
rect 10284 16136 10692 16164
rect 10284 16124 10290 16136
rect 10686 16124 10692 16136
rect 10744 16124 10750 16176
rect 11808 16164 11836 16204
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 13722 16232 13728 16244
rect 11931 16204 13728 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 15378 16192 15384 16244
rect 15436 16232 15442 16244
rect 16025 16235 16083 16241
rect 16025 16232 16037 16235
rect 15436 16204 16037 16232
rect 15436 16192 15442 16204
rect 16025 16201 16037 16204
rect 16071 16201 16083 16235
rect 16942 16232 16948 16244
rect 16903 16204 16948 16232
rect 16025 16195 16083 16201
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 19886 16232 19892 16244
rect 17276 16204 19892 16232
rect 17276 16192 17282 16204
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 20530 16192 20536 16244
rect 20588 16232 20594 16244
rect 22005 16235 22063 16241
rect 22005 16232 22017 16235
rect 20588 16204 22017 16232
rect 20588 16192 20594 16204
rect 22005 16201 22017 16204
rect 22051 16201 22063 16235
rect 22005 16195 22063 16201
rect 12529 16167 12587 16173
rect 11808 16136 12480 16164
rect 5534 16096 5540 16108
rect 5276 16068 5540 16096
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 5905 16099 5963 16105
rect 5905 16096 5917 16099
rect 5776 16068 5917 16096
rect 5776 16056 5782 16068
rect 5905 16065 5917 16068
rect 5951 16065 5963 16099
rect 5905 16059 5963 16065
rect 5997 16099 6055 16105
rect 5997 16065 6009 16099
rect 6043 16096 6055 16099
rect 6917 16099 6975 16105
rect 6917 16096 6929 16099
rect 6043 16068 6929 16096
rect 6043 16065 6055 16068
rect 5997 16059 6055 16065
rect 6917 16065 6929 16068
rect 6963 16096 6975 16099
rect 7006 16096 7012 16108
rect 6963 16068 7012 16096
rect 6963 16065 6975 16068
rect 6917 16059 6975 16065
rect 7006 16056 7012 16068
rect 7064 16056 7070 16108
rect 7392 16096 7420 16124
rect 7116 16068 7420 16096
rect 9401 16099 9459 16105
rect 4522 15988 4528 16040
rect 4580 16028 4586 16040
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 4580 16000 4629 16028
rect 4580 15988 4586 16000
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 5166 15988 5172 16040
rect 5224 16028 5230 16040
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 5224 16000 6837 16028
rect 5224 15988 5230 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 7116 16028 7144 16068
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 10778 16096 10784 16108
rect 9447 16068 10784 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10962 16096 10968 16108
rect 10923 16068 10968 16096
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 12452 16105 12480 16136
rect 12529 16133 12541 16167
rect 12575 16164 12587 16167
rect 13265 16167 13323 16173
rect 13265 16164 13277 16167
rect 12575 16136 13277 16164
rect 12575 16133 12587 16136
rect 12529 16127 12587 16133
rect 13265 16133 13277 16136
rect 13311 16133 13323 16167
rect 13265 16127 13323 16133
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 14461 16167 14519 16173
rect 14461 16164 14473 16167
rect 14424 16136 14473 16164
rect 14424 16124 14430 16136
rect 14461 16133 14473 16136
rect 14507 16133 14519 16167
rect 14461 16127 14519 16133
rect 17310 16124 17316 16176
rect 17368 16164 17374 16176
rect 18509 16167 18567 16173
rect 18509 16164 18521 16167
rect 17368 16136 18521 16164
rect 17368 16124 17374 16136
rect 18509 16133 18521 16136
rect 18555 16133 18567 16167
rect 18509 16127 18567 16133
rect 19334 16124 19340 16176
rect 19392 16164 19398 16176
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 19392 16136 19717 16164
rect 19392 16124 19398 16136
rect 19705 16133 19717 16136
rect 19751 16133 19763 16167
rect 19705 16127 19763 16133
rect 19794 16124 19800 16176
rect 19852 16164 19858 16176
rect 20349 16167 20407 16173
rect 20349 16164 20361 16167
rect 19852 16136 20361 16164
rect 19852 16124 19858 16136
rect 20349 16133 20361 16136
rect 20395 16133 20407 16167
rect 20349 16127 20407 16133
rect 11793 16099 11851 16105
rect 11793 16065 11805 16099
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16096 12495 16099
rect 16114 16096 16120 16108
rect 12483 16068 12940 16096
rect 16075 16068 16120 16096
rect 12483 16065 12495 16068
rect 12437 16059 12495 16065
rect 6825 15991 6883 15997
rect 6932 16000 7144 16028
rect 7377 16031 7435 16037
rect 1673 15963 1731 15969
rect 1673 15929 1685 15963
rect 1719 15960 1731 15963
rect 2774 15960 2780 15972
rect 1719 15932 2780 15960
rect 1719 15929 1731 15932
rect 1673 15923 1731 15929
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 5258 15920 5264 15972
rect 5316 15960 5322 15972
rect 6932 15960 6960 16000
rect 7377 15997 7389 16031
rect 7423 15997 7435 16031
rect 11808 16028 11836 16059
rect 10244 16016 11836 16028
rect 7377 15991 7435 15997
rect 10060 16000 11836 16016
rect 5316 15932 6960 15960
rect 5316 15920 5322 15932
rect 7006 15920 7012 15972
rect 7064 15960 7070 15972
rect 7282 15960 7288 15972
rect 7064 15932 7288 15960
rect 7064 15920 7070 15932
rect 7282 15920 7288 15932
rect 7340 15960 7346 15972
rect 7392 15960 7420 15991
rect 10060 15988 10272 16000
rect 10060 15960 10088 15988
rect 10318 15960 10324 15972
rect 7340 15932 7420 15960
rect 8680 15932 10088 15960
rect 10279 15932 10324 15960
rect 7340 15920 7346 15932
rect 2314 15892 2320 15904
rect 2275 15864 2320 15892
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 2498 15852 2504 15904
rect 2556 15892 2562 15904
rect 8680 15892 8708 15932
rect 10318 15920 10324 15932
rect 10376 15920 10382 15972
rect 2556 15864 8708 15892
rect 11057 15895 11115 15901
rect 2556 15852 2562 15864
rect 11057 15861 11069 15895
rect 11103 15892 11115 15895
rect 12802 15892 12808 15904
rect 11103 15864 12808 15892
rect 11103 15861 11115 15864
rect 11057 15855 11115 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 12912 15892 12940 16068
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16850 16096 16856 16108
rect 16811 16068 16856 16096
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 22554 16096 22560 16108
rect 22515 16068 22560 16096
rect 22554 16056 22560 16068
rect 22612 16056 22618 16108
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 35713 16099 35771 16105
rect 35713 16065 35725 16099
rect 35759 16096 35771 16099
rect 36354 16096 36360 16108
rect 35759 16068 36360 16096
rect 35759 16065 35771 16068
rect 35713 16059 35771 16065
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 13173 16031 13231 16037
rect 13044 16016 13124 16028
rect 13173 16016 13185 16031
rect 13044 16000 13185 16016
rect 13044 15988 13050 16000
rect 13096 15997 13185 16000
rect 13219 15997 13231 16031
rect 13096 15991 13231 15997
rect 13096 15988 13205 15991
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14369 16031 14427 16037
rect 14369 16028 14381 16031
rect 14148 16000 14381 16028
rect 14148 15988 14154 16000
rect 14369 15997 14381 16000
rect 14415 16028 14427 16031
rect 14918 16028 14924 16040
rect 14415 16000 14924 16028
rect 14415 15997 14427 16000
rect 14369 15991 14427 15997
rect 14918 15988 14924 16000
rect 14976 15988 14982 16040
rect 15286 16028 15292 16040
rect 15247 16000 15292 16028
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 16206 15988 16212 16040
rect 16264 16028 16270 16040
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 16264 16000 17969 16028
rect 16264 15988 16270 16000
rect 17957 15997 17969 16000
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 18601 16031 18659 16037
rect 18601 15997 18613 16031
rect 18647 16028 18659 16031
rect 19797 16031 19855 16037
rect 18647 16000 19380 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 13725 15963 13783 15969
rect 13725 15929 13737 15963
rect 13771 15960 13783 15963
rect 16574 15960 16580 15972
rect 13771 15932 16580 15960
rect 13771 15929 13783 15932
rect 13725 15923 13783 15929
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 17972 15960 18000 15991
rect 19245 15963 19303 15969
rect 19245 15960 19257 15963
rect 17972 15932 19257 15960
rect 19245 15929 19257 15932
rect 19291 15929 19303 15963
rect 19352 15960 19380 16000
rect 19797 15997 19809 16031
rect 19843 16028 19855 16031
rect 20070 16028 20076 16040
rect 19843 16000 20076 16028
rect 19843 15997 19855 16000
rect 19797 15991 19855 15997
rect 20070 15988 20076 16000
rect 20128 15988 20134 16040
rect 20622 15988 20628 16040
rect 20680 16028 20686 16040
rect 26329 16031 26387 16037
rect 26329 16028 26341 16031
rect 20680 16000 26341 16028
rect 20680 15988 20686 16000
rect 26329 15997 26341 16000
rect 26375 15997 26387 16031
rect 26329 15991 26387 15997
rect 20162 15960 20168 15972
rect 19352 15932 20168 15960
rect 19245 15923 19303 15929
rect 20162 15920 20168 15932
rect 20220 15920 20226 15972
rect 16022 15892 16028 15904
rect 12912 15864 16028 15892
rect 16022 15852 16028 15864
rect 16080 15892 16086 15904
rect 17494 15892 17500 15904
rect 16080 15864 17500 15892
rect 16080 15852 16086 15864
rect 17494 15852 17500 15864
rect 17552 15892 17558 15904
rect 18506 15892 18512 15904
rect 17552 15864 18512 15892
rect 17552 15852 17558 15864
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 18782 15852 18788 15904
rect 18840 15892 18846 15904
rect 20993 15895 21051 15901
rect 20993 15892 21005 15895
rect 18840 15864 21005 15892
rect 18840 15852 18846 15864
rect 20993 15861 21005 15864
rect 21039 15861 21051 15895
rect 26436 15892 26464 16059
rect 36354 16056 36360 16068
rect 36412 16056 36418 16108
rect 35894 15892 35900 15904
rect 26436 15864 35900 15892
rect 20993 15855 21051 15861
rect 35894 15852 35900 15864
rect 35952 15892 35958 15904
rect 36173 15895 36231 15901
rect 36173 15892 36185 15895
rect 35952 15864 36185 15892
rect 35952 15852 35958 15864
rect 36173 15861 36185 15864
rect 36219 15861 36231 15895
rect 36173 15855 36231 15861
rect 1104 15802 36892 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 36892 15802
rect 1104 15728 36892 15750
rect 3329 15691 3387 15697
rect 3329 15657 3341 15691
rect 3375 15688 3387 15691
rect 6454 15688 6460 15700
rect 3375 15660 6460 15688
rect 3375 15657 3387 15660
rect 3329 15651 3387 15657
rect 6454 15648 6460 15660
rect 6512 15648 6518 15700
rect 8570 15688 8576 15700
rect 6564 15660 8576 15688
rect 1578 15552 1584 15564
rect 1539 15524 1584 15552
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 6564 15552 6592 15660
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 8938 15648 8944 15700
rect 8996 15688 9002 15700
rect 10870 15688 10876 15700
rect 8996 15660 10876 15688
rect 8996 15648 9002 15660
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 14458 15688 14464 15700
rect 12406 15660 14464 15688
rect 2976 15524 6592 15552
rect 8297 15555 8355 15561
rect 2976 15470 3004 15524
rect 8297 15521 8309 15555
rect 8343 15552 8355 15555
rect 8662 15552 8668 15564
rect 8343 15524 8668 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 8662 15512 8668 15524
rect 8720 15552 8726 15564
rect 12406 15552 12434 15660
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 17310 15688 17316 15700
rect 17271 15660 17316 15688
rect 17310 15648 17316 15660
rect 17368 15648 17374 15700
rect 18690 15688 18696 15700
rect 18651 15660 18696 15688
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 21637 15691 21695 15697
rect 21637 15688 21649 15691
rect 18800 15660 21649 15688
rect 18800 15620 18828 15660
rect 21637 15657 21649 15660
rect 21683 15657 21695 15691
rect 21637 15651 21695 15657
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 30558 15688 30564 15700
rect 22612 15660 30564 15688
rect 22612 15648 22618 15660
rect 30558 15648 30564 15660
rect 30616 15648 30622 15700
rect 14752 15592 18828 15620
rect 8720 15524 12434 15552
rect 12529 15555 12587 15561
rect 8720 15512 8726 15524
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 13725 15555 13783 15561
rect 13725 15552 13737 15555
rect 12575 15524 13737 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 13725 15521 13737 15524
rect 13771 15552 13783 15555
rect 14182 15552 14188 15564
rect 13771 15524 14188 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4212 15456 4261 15484
rect 4212 15444 4218 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 6362 15444 6368 15496
rect 6420 15484 6426 15496
rect 6549 15487 6607 15493
rect 6549 15484 6561 15487
rect 6420 15456 6561 15484
rect 6420 15444 6426 15456
rect 6549 15453 6561 15456
rect 6595 15453 6607 15487
rect 6549 15447 6607 15453
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8628 15456 9137 15484
rect 8628 15444 8634 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 14090 15444 14096 15496
rect 14148 15484 14154 15496
rect 14752 15493 14780 15592
rect 19886 15580 19892 15632
rect 19944 15620 19950 15632
rect 19981 15623 20039 15629
rect 19981 15620 19993 15623
rect 19944 15592 19993 15620
rect 19944 15580 19950 15592
rect 19981 15589 19993 15592
rect 20027 15589 20039 15623
rect 19981 15583 20039 15589
rect 20622 15580 20628 15632
rect 20680 15580 20686 15632
rect 15473 15555 15531 15561
rect 15473 15521 15485 15555
rect 15519 15552 15531 15555
rect 15562 15552 15568 15564
rect 15519 15524 15568 15552
rect 15519 15521 15531 15524
rect 15473 15515 15531 15521
rect 15562 15512 15568 15524
rect 15620 15552 15626 15564
rect 16298 15552 16304 15564
rect 15620 15524 16304 15552
rect 15620 15512 15626 15524
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 20254 15552 20260 15564
rect 17144 15524 20260 15552
rect 14737 15487 14795 15493
rect 14737 15484 14749 15487
rect 14148 15456 14749 15484
rect 14148 15444 14154 15456
rect 14737 15453 14749 15456
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 16117 15487 16175 15493
rect 16117 15453 16129 15487
rect 16163 15484 16175 15487
rect 17144 15484 17172 15524
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 20640 15552 20668 15580
rect 20579 15524 20668 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 16163 15456 17172 15484
rect 17221 15487 17279 15493
rect 16163 15453 16175 15456
rect 16117 15447 16175 15453
rect 17221 15453 17233 15487
rect 17267 15484 17279 15487
rect 17310 15484 17316 15496
rect 17267 15456 17316 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 1394 15376 1400 15428
rect 1452 15416 1458 15428
rect 1857 15419 1915 15425
rect 1857 15416 1869 15419
rect 1452 15388 1869 15416
rect 1452 15376 1458 15388
rect 1857 15385 1869 15388
rect 1903 15385 1915 15419
rect 1857 15379 1915 15385
rect 4525 15419 4583 15425
rect 4525 15385 4537 15419
rect 4571 15416 4583 15419
rect 6086 15416 6092 15428
rect 4571 15388 4752 15416
rect 5750 15388 6092 15416
rect 4571 15385 4583 15388
rect 4525 15379 4583 15385
rect 4724 15360 4752 15388
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 9401 15419 9459 15425
rect 7866 15388 8248 15416
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 4890 15348 4896 15360
rect 4764 15320 4896 15348
rect 4764 15308 4770 15320
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 5997 15351 6055 15357
rect 5997 15317 6009 15351
rect 6043 15348 6055 15351
rect 7374 15348 7380 15360
rect 6043 15320 7380 15348
rect 6043 15317 6055 15320
rect 5997 15311 6055 15317
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 8220 15348 8248 15388
rect 9401 15385 9413 15419
rect 9447 15416 9459 15419
rect 9490 15416 9496 15428
rect 9447 15388 9496 15416
rect 9447 15385 9459 15388
rect 9401 15379 9459 15385
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 11885 15419 11943 15425
rect 11885 15416 11897 15419
rect 11112 15388 11897 15416
rect 11112 15376 11118 15388
rect 11885 15385 11897 15388
rect 11931 15385 11943 15419
rect 11885 15379 11943 15385
rect 11977 15419 12035 15425
rect 11977 15385 11989 15419
rect 12023 15416 12035 15419
rect 12023 15388 12434 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 10042 15348 10048 15360
rect 8220 15320 10048 15348
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 11900 15348 11928 15379
rect 12158 15348 12164 15360
rect 11900 15320 12164 15348
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 12406 15348 12434 15388
rect 12802 15376 12808 15428
rect 12860 15416 12866 15428
rect 13078 15416 13084 15428
rect 12860 15388 13084 15416
rect 12860 15376 12866 15388
rect 13078 15376 13084 15388
rect 13136 15376 13142 15428
rect 13173 15419 13231 15425
rect 13173 15385 13185 15419
rect 13219 15385 13231 15419
rect 15286 15416 15292 15428
rect 13173 15379 13231 15385
rect 14752 15388 15292 15416
rect 12986 15348 12992 15360
rect 12406 15320 12992 15348
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 13188 15348 13216 15379
rect 14752 15348 14780 15388
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 15565 15419 15623 15425
rect 15565 15385 15577 15419
rect 15611 15385 15623 15419
rect 15565 15379 15623 15385
rect 13188 15320 14780 15348
rect 14829 15351 14887 15357
rect 14829 15317 14841 15351
rect 14875 15348 14887 15351
rect 15580 15348 15608 15379
rect 15746 15376 15752 15428
rect 15804 15416 15810 15428
rect 16132 15416 16160 15447
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15484 18107 15487
rect 18138 15484 18144 15496
rect 18095 15456 18144 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15486 18659 15487
rect 18647 15458 18736 15486
rect 18647 15453 18659 15458
rect 18601 15447 18659 15453
rect 15804 15388 16160 15416
rect 17328 15416 17356 15444
rect 17586 15416 17592 15428
rect 17328 15388 17592 15416
rect 15804 15376 15810 15388
rect 17586 15376 17592 15388
rect 17644 15416 17650 15428
rect 18708 15416 18736 15458
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 19794 15484 19800 15496
rect 19024 15456 19800 15484
rect 19024 15444 19030 15456
rect 19794 15444 19800 15456
rect 19852 15444 19858 15496
rect 20898 15444 20904 15496
rect 20956 15484 20962 15496
rect 22741 15487 22799 15493
rect 22741 15484 22753 15487
rect 20956 15456 22753 15484
rect 20956 15444 20962 15456
rect 22741 15453 22753 15456
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 18782 15416 18788 15428
rect 17644 15388 18276 15416
rect 18708 15388 18788 15416
rect 17644 15376 17650 15388
rect 16758 15348 16764 15360
rect 14875 15320 15608 15348
rect 16719 15320 16764 15348
rect 14875 15317 14887 15320
rect 14829 15311 14887 15317
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 17770 15308 17776 15360
rect 17828 15348 17834 15360
rect 17957 15351 18015 15357
rect 17957 15348 17969 15351
rect 17828 15320 17969 15348
rect 17828 15308 17834 15320
rect 17957 15317 17969 15320
rect 18003 15317 18015 15351
rect 18248 15348 18276 15388
rect 18782 15376 18788 15388
rect 18840 15376 18846 15428
rect 20438 15416 20444 15428
rect 20399 15388 20444 15416
rect 20438 15376 20444 15388
rect 20496 15376 20502 15428
rect 22186 15416 22192 15428
rect 22147 15388 22192 15416
rect 22186 15376 22192 15388
rect 22244 15376 22250 15428
rect 21085 15351 21143 15357
rect 21085 15348 21097 15351
rect 18248 15320 21097 15348
rect 17957 15311 18015 15317
rect 21085 15317 21097 15320
rect 21131 15317 21143 15351
rect 21085 15311 21143 15317
rect 1104 15258 36892 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 36892 15258
rect 1104 15184 36892 15206
rect 3050 15144 3056 15156
rect 1596 15116 3056 15144
rect 1596 15085 1624 15116
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 5537 15147 5595 15153
rect 5537 15144 5549 15147
rect 5408 15116 5549 15144
rect 5408 15104 5414 15116
rect 5537 15113 5549 15116
rect 5583 15113 5595 15147
rect 10318 15144 10324 15156
rect 5537 15107 5595 15113
rect 6748 15116 10324 15144
rect 1581 15079 1639 15085
rect 1581 15045 1593 15079
rect 1627 15045 1639 15079
rect 1581 15039 1639 15045
rect 2866 15036 2872 15088
rect 2924 15036 2930 15088
rect 3329 15079 3387 15085
rect 3329 15045 3341 15079
rect 3375 15076 3387 15079
rect 3418 15076 3424 15088
rect 3375 15048 3424 15076
rect 3375 15045 3387 15048
rect 3329 15039 3387 15045
rect 3418 15036 3424 15048
rect 3476 15036 3482 15088
rect 3786 15036 3792 15088
rect 3844 15076 3850 15088
rect 6641 15079 6699 15085
rect 6641 15076 6653 15079
rect 3844 15048 6653 15076
rect 3844 15036 3850 15048
rect 6641 15045 6653 15048
rect 6687 15045 6699 15079
rect 6641 15039 6699 15045
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 6748 15017 6776 15116
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 11054 15144 11060 15156
rect 10796 15116 11060 15144
rect 10796 15076 10824 15116
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 11793 15147 11851 15153
rect 11793 15113 11805 15147
rect 11839 15144 11851 15147
rect 11882 15144 11888 15156
rect 11839 15116 11888 15144
rect 11839 15113 11851 15116
rect 11793 15107 11851 15113
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 13446 15144 13452 15156
rect 13320 15116 13452 15144
rect 13320 15104 13326 15116
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 15102 15144 15108 15156
rect 14108 15116 15108 15144
rect 10962 15076 10968 15088
rect 8786 15048 10824 15076
rect 10923 15048 10968 15076
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11330 15036 11336 15088
rect 11388 15076 11394 15088
rect 12805 15079 12863 15085
rect 12805 15076 12817 15079
rect 11388 15048 12817 15076
rect 11388 15036 11394 15048
rect 12805 15045 12817 15048
rect 12851 15045 12863 15079
rect 12805 15039 12863 15045
rect 13357 15079 13415 15085
rect 13357 15045 13369 15079
rect 13403 15076 13415 15079
rect 13630 15076 13636 15088
rect 13403 15048 13636 15076
rect 13403 15045 13415 15048
rect 13357 15039 13415 15045
rect 13630 15036 13636 15048
rect 13688 15036 13694 15088
rect 14108 15076 14136 15116
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 17862 15144 17868 15156
rect 15212 15116 17868 15144
rect 13924 15048 14136 15076
rect 14185 15079 14243 15085
rect 4249 15011 4307 15017
rect 4249 15008 4261 15011
rect 4120 14980 4261 15008
rect 4120 14968 4126 14980
rect 4249 14977 4261 14980
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 9953 15011 10011 15017
rect 9953 14977 9965 15011
rect 9999 15008 10011 15011
rect 10410 15008 10416 15020
rect 9999 14980 10416 15008
rect 9999 14977 10011 14980
rect 9953 14971 10011 14977
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 11701 15011 11759 15017
rect 11296 14980 11652 15008
rect 11296 14968 11302 14980
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14940 3663 14943
rect 3970 14940 3976 14952
rect 3651 14912 3976 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 3970 14900 3976 14912
rect 4028 14940 4034 14952
rect 4154 14940 4160 14952
rect 4028 14912 4160 14940
rect 4028 14900 4034 14912
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 6972 14912 7297 14940
rect 6972 14900 6978 14912
rect 7285 14909 7297 14912
rect 7331 14909 7343 14943
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7285 14903 7343 14909
rect 7392 14912 7573 14940
rect 3878 14832 3884 14884
rect 3936 14872 3942 14884
rect 7392 14872 7420 14912
rect 7561 14909 7573 14912
rect 7607 14909 7619 14943
rect 7561 14903 7619 14909
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 8352 14912 9321 14940
rect 8352 14900 8358 14912
rect 9309 14909 9321 14912
rect 9355 14940 9367 14943
rect 9398 14940 9404 14952
rect 9355 14912 9404 14940
rect 9355 14909 9367 14912
rect 9309 14903 9367 14909
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 10686 14940 10692 14952
rect 10647 14912 10692 14940
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 11057 14943 11115 14949
rect 11057 14909 11069 14943
rect 11103 14940 11115 14943
rect 11330 14940 11336 14952
rect 11103 14912 11336 14940
rect 11103 14909 11115 14912
rect 11057 14903 11115 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 11624 14940 11652 14980
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 11790 15008 11796 15020
rect 11747 14980 11796 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 13449 14943 13507 14949
rect 11624 14912 13400 14940
rect 3936 14844 7420 14872
rect 3936 14832 3942 14844
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 13262 14872 13268 14884
rect 12584 14844 13268 14872
rect 12584 14832 12590 14844
rect 13262 14832 13268 14844
rect 13320 14832 13326 14884
rect 13372 14872 13400 14912
rect 13449 14909 13461 14943
rect 13495 14940 13507 14943
rect 13924 14940 13952 15048
rect 14185 15045 14197 15079
rect 14231 15076 14243 15079
rect 15010 15076 15016 15088
rect 14231 15048 15016 15076
rect 14231 15045 14243 15048
rect 14185 15039 14243 15045
rect 15010 15036 15016 15048
rect 15068 15036 15074 15088
rect 15212 15076 15240 15116
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 18141 15147 18199 15153
rect 18141 15113 18153 15147
rect 18187 15144 18199 15147
rect 20438 15144 20444 15156
rect 18187 15116 20444 15144
rect 18187 15113 18199 15116
rect 18141 15107 18199 15113
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 15378 15076 15384 15088
rect 15120 15048 15240 15076
rect 15339 15048 15384 15076
rect 14737 15011 14795 15017
rect 14737 14977 14749 15011
rect 14783 15008 14795 15011
rect 15120 15008 15148 15048
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 16945 15079 17003 15085
rect 16945 15076 16957 15079
rect 16816 15048 16957 15076
rect 16816 15036 16822 15048
rect 16945 15045 16957 15048
rect 16991 15045 17003 15079
rect 16945 15039 17003 15045
rect 17037 15079 17095 15085
rect 17037 15045 17049 15079
rect 17083 15076 17095 15079
rect 17954 15076 17960 15088
rect 17083 15048 17960 15076
rect 17083 15045 17095 15048
rect 17037 15039 17095 15045
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 18598 15036 18604 15088
rect 18656 15076 18662 15088
rect 18693 15079 18751 15085
rect 18693 15076 18705 15079
rect 18656 15048 18705 15076
rect 18656 15036 18662 15048
rect 18693 15045 18705 15048
rect 18739 15045 18751 15079
rect 18693 15039 18751 15045
rect 19337 15079 19395 15085
rect 19337 15045 19349 15079
rect 19383 15076 19395 15079
rect 20073 15079 20131 15085
rect 20073 15076 20085 15079
rect 19383 15048 20085 15076
rect 19383 15045 19395 15048
rect 19337 15039 19395 15045
rect 20073 15045 20085 15048
rect 20119 15045 20131 15079
rect 20073 15039 20131 15045
rect 14783 14980 15148 15008
rect 14783 14977 14795 14980
rect 14737 14971 14795 14977
rect 17586 14968 17592 15020
rect 17644 15008 17650 15020
rect 18049 15011 18107 15017
rect 18049 15008 18061 15011
rect 17644 14980 18061 15008
rect 17644 14968 17650 14980
rect 18049 14977 18061 14980
rect 18095 15008 18107 15011
rect 18322 15008 18328 15020
rect 18095 14980 18328 15008
rect 18095 14977 18107 14980
rect 18049 14971 18107 14977
rect 18322 14968 18328 14980
rect 18380 14968 18386 15020
rect 18708 15008 18736 15039
rect 20254 15036 20260 15088
rect 20312 15076 20318 15088
rect 20625 15079 20683 15085
rect 20625 15076 20637 15079
rect 20312 15048 20637 15076
rect 20312 15036 20318 15048
rect 20625 15045 20637 15048
rect 20671 15076 20683 15079
rect 21174 15076 21180 15088
rect 20671 15048 21180 15076
rect 20671 15045 20683 15048
rect 20625 15039 20683 15045
rect 21174 15036 21180 15048
rect 21232 15036 21238 15088
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 18708 14980 19257 15008
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 20772 14980 21097 15008
rect 20772 14968 20778 14980
rect 21085 14977 21097 14980
rect 21131 15008 21143 15011
rect 21266 15008 21272 15020
rect 21131 14980 21272 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 13495 14912 13952 14940
rect 14093 14943 14151 14949
rect 13495 14909 13507 14912
rect 13449 14903 13507 14909
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14182 14940 14188 14952
rect 14139 14912 14188 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 15289 14943 15347 14949
rect 15289 14940 15301 14943
rect 14516 14912 15301 14940
rect 14516 14900 14522 14912
rect 15289 14909 15301 14912
rect 15335 14909 15347 14943
rect 15654 14940 15660 14952
rect 15615 14912 15660 14940
rect 15289 14903 15347 14909
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 17218 14940 17224 14952
rect 17179 14912 17224 14940
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14940 20039 14943
rect 20070 14940 20076 14952
rect 20027 14912 20076 14940
rect 20027 14909 20039 14912
rect 19981 14903 20039 14909
rect 20070 14900 20076 14912
rect 20128 14940 20134 14952
rect 20622 14940 20628 14952
rect 20128 14912 20628 14940
rect 20128 14900 20134 14912
rect 20622 14900 20628 14912
rect 20680 14940 20686 14952
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 20680 14912 21189 14940
rect 20680 14900 20686 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 22557 14943 22615 14949
rect 22557 14940 22569 14943
rect 21177 14903 21235 14909
rect 22066 14912 22569 14940
rect 13814 14872 13820 14884
rect 13372 14844 13820 14872
rect 13814 14832 13820 14844
rect 13872 14832 13878 14884
rect 22066 14872 22094 14912
rect 22557 14909 22569 14912
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 17236 14844 22094 14872
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 2648 14776 9873 14804
rect 2648 14764 2654 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 9861 14767 9919 14773
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 17236 14804 17264 14844
rect 11848 14776 17264 14804
rect 11848 14764 11854 14776
rect 21266 14764 21272 14816
rect 21324 14804 21330 14816
rect 22097 14807 22155 14813
rect 22097 14804 22109 14807
rect 21324 14776 22109 14804
rect 21324 14764 21330 14776
rect 22097 14773 22109 14776
rect 22143 14804 22155 14807
rect 23474 14804 23480 14816
rect 22143 14776 23480 14804
rect 22143 14773 22155 14776
rect 22097 14767 22155 14773
rect 23474 14764 23480 14776
rect 23532 14764 23538 14816
rect 1104 14714 36892 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 36892 14714
rect 1104 14640 36892 14662
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 3602 14600 3608 14612
rect 3467 14572 3608 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 4801 14603 4859 14609
rect 4801 14569 4813 14603
rect 4847 14600 4859 14603
rect 7006 14600 7012 14612
rect 4847 14572 7012 14600
rect 4847 14569 4859 14572
rect 4801 14563 4859 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7300 14572 8524 14600
rect 2958 14492 2964 14544
rect 3016 14532 3022 14544
rect 5718 14532 5724 14544
rect 3016 14504 5724 14532
rect 3016 14492 3022 14504
rect 5718 14492 5724 14504
rect 5776 14492 5782 14544
rect 6178 14492 6184 14544
rect 6236 14532 6242 14544
rect 7300 14532 7328 14572
rect 6236 14504 7328 14532
rect 8496 14532 8524 14572
rect 9398 14560 9404 14612
rect 9456 14600 9462 14612
rect 12526 14600 12532 14612
rect 9456 14572 12532 14600
rect 9456 14560 9462 14572
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 12986 14600 12992 14612
rect 12947 14572 12992 14600
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 13630 14600 13636 14612
rect 13591 14572 13636 14600
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 15010 14600 15016 14612
rect 14971 14572 15016 14600
rect 15010 14560 15016 14572
rect 15068 14560 15074 14612
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 16025 14603 16083 14609
rect 16025 14600 16037 14603
rect 15344 14572 16037 14600
rect 15344 14560 15350 14572
rect 16025 14569 16037 14572
rect 16071 14569 16083 14603
rect 16025 14563 16083 14569
rect 16114 14560 16120 14612
rect 16172 14600 16178 14612
rect 18782 14600 18788 14612
rect 16172 14572 18788 14600
rect 16172 14560 16178 14572
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 22186 14532 22192 14544
rect 8496 14504 9260 14532
rect 6236 14492 6242 14504
rect 1578 14424 1584 14476
rect 1636 14464 1642 14476
rect 1673 14467 1731 14473
rect 1673 14464 1685 14467
rect 1636 14436 1685 14464
rect 1636 14424 1642 14436
rect 1673 14433 1685 14436
rect 1719 14433 1731 14467
rect 1673 14427 1731 14433
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2038 14464 2044 14476
rect 1995 14436 2044 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 2406 14424 2412 14476
rect 2464 14464 2470 14476
rect 6822 14464 6828 14476
rect 2464 14436 6828 14464
rect 2464 14424 2470 14436
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 8570 14464 8576 14476
rect 6972 14436 8576 14464
rect 6972 14424 6978 14436
rect 8570 14424 8576 14436
rect 8628 14464 8634 14476
rect 9125 14467 9183 14473
rect 9125 14464 9137 14467
rect 8628 14436 9137 14464
rect 8628 14424 8634 14436
rect 9125 14433 9137 14436
rect 9171 14433 9183 14467
rect 9232 14464 9260 14504
rect 10428 14504 20116 14532
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 9232 14436 9413 14464
rect 9125 14427 9183 14433
rect 9401 14433 9413 14436
rect 9447 14464 9459 14467
rect 10428 14464 10456 14504
rect 9447 14436 10456 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 12342 14424 12348 14476
rect 12400 14464 12406 14476
rect 18046 14464 18052 14476
rect 12400 14436 15148 14464
rect 18007 14436 18052 14464
rect 12400 14424 12406 14436
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 6089 14399 6147 14405
rect 6089 14396 6101 14399
rect 5408 14368 6101 14396
rect 5408 14356 5414 14368
rect 6089 14365 6101 14368
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 13081 14399 13139 14405
rect 10836 14368 11468 14396
rect 10836 14356 10842 14368
rect 5258 14328 5264 14340
rect 3174 14300 5264 14328
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 6549 14331 6607 14337
rect 6549 14297 6561 14331
rect 6595 14328 6607 14331
rect 7006 14328 7012 14340
rect 6595 14300 7012 14328
rect 6595 14297 6607 14300
rect 6549 14291 6607 14297
rect 7006 14288 7012 14300
rect 7064 14288 7070 14340
rect 7834 14288 7840 14340
rect 7892 14288 7898 14340
rect 8294 14328 8300 14340
rect 8207 14300 8300 14328
rect 8294 14288 8300 14300
rect 8352 14328 8358 14340
rect 8754 14328 8760 14340
rect 8352 14300 8760 14328
rect 8352 14288 8358 14300
rect 8754 14288 8760 14300
rect 8812 14288 8818 14340
rect 11440 14337 11468 14368
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13354 14396 13360 14408
rect 13127 14368 13360 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 13538 14356 13544 14408
rect 13596 14396 13602 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13596 14368 13737 14396
rect 13596 14356 13602 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 14458 14396 14464 14408
rect 14419 14368 14464 14396
rect 13725 14359 13783 14365
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 15120 14405 15148 14436
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 19978 14464 19984 14476
rect 19939 14436 19984 14464
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 20088 14464 20116 14504
rect 20364 14504 22192 14532
rect 20364 14464 20392 14504
rect 22186 14492 22192 14504
rect 22244 14492 22250 14544
rect 20088 14436 20392 14464
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 20680 14436 22385 14464
rect 20680 14424 20686 14436
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 22373 14427 22431 14433
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14396 16175 14399
rect 16390 14396 16396 14408
rect 16163 14368 16396 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 11425 14331 11483 14337
rect 9416 14300 9890 14328
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 4522 14260 4528 14272
rect 3568 14232 4528 14260
rect 3568 14220 3574 14232
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 9416 14260 9444 14300
rect 11425 14297 11437 14331
rect 11471 14297 11483 14331
rect 11974 14328 11980 14340
rect 11935 14300 11980 14328
rect 11425 14291 11483 14297
rect 11974 14288 11980 14300
rect 12032 14288 12038 14340
rect 12066 14288 12072 14340
rect 12124 14328 12130 14340
rect 16132 14328 16160 14359
rect 16390 14356 16396 14368
rect 16448 14356 16454 14408
rect 36081 14399 36139 14405
rect 36081 14396 36093 14399
rect 35866 14368 36093 14396
rect 12124 14300 12169 14328
rect 15120 14300 16160 14328
rect 17129 14331 17187 14337
rect 12124 14288 12130 14300
rect 5868 14232 9444 14260
rect 5868 14220 5874 14232
rect 9582 14220 9588 14272
rect 9640 14260 9646 14272
rect 10134 14260 10140 14272
rect 9640 14232 10140 14260
rect 9640 14220 9646 14232
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 10873 14263 10931 14269
rect 10873 14260 10885 14263
rect 10836 14232 10885 14260
rect 10836 14220 10842 14232
rect 10873 14229 10885 14232
rect 10919 14229 10931 14263
rect 10873 14223 10931 14229
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 15120 14260 15148 14300
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 17681 14331 17739 14337
rect 17681 14328 17693 14331
rect 17175 14300 17693 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 17681 14297 17693 14300
rect 17727 14297 17739 14331
rect 17681 14291 17739 14297
rect 17773 14331 17831 14337
rect 17773 14297 17785 14331
rect 17819 14297 17831 14331
rect 17773 14291 17831 14297
rect 13688 14232 15148 14260
rect 13688 14220 13694 14232
rect 15286 14220 15292 14272
rect 15344 14260 15350 14272
rect 17788 14260 17816 14291
rect 20070 14288 20076 14340
rect 20128 14328 20134 14340
rect 20625 14331 20683 14337
rect 20128 14300 20173 14328
rect 20128 14288 20134 14300
rect 20625 14297 20637 14331
rect 20671 14297 20683 14331
rect 21082 14328 21088 14340
rect 21043 14300 21088 14328
rect 20625 14291 20683 14297
rect 15344 14232 17816 14260
rect 15344 14220 15350 14232
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 20640 14260 20668 14291
rect 21082 14288 21088 14300
rect 21140 14288 21146 14340
rect 21634 14328 21640 14340
rect 21595 14300 21640 14328
rect 21634 14288 21640 14300
rect 21692 14288 21698 14340
rect 21726 14288 21732 14340
rect 21784 14328 21790 14340
rect 21784 14300 21829 14328
rect 21784 14288 21790 14300
rect 22462 14288 22468 14340
rect 22520 14328 22526 14340
rect 23017 14331 23075 14337
rect 22520 14300 22565 14328
rect 22520 14288 22526 14300
rect 23017 14297 23029 14331
rect 23063 14297 23075 14331
rect 23017 14291 23075 14297
rect 22738 14260 22744 14272
rect 17920 14232 22744 14260
rect 17920 14220 17926 14232
rect 22738 14220 22744 14232
rect 22796 14260 22802 14272
rect 23032 14260 23060 14291
rect 35526 14260 35532 14272
rect 22796 14232 23060 14260
rect 35487 14232 35532 14260
rect 22796 14220 22802 14232
rect 35526 14220 35532 14232
rect 35584 14260 35590 14272
rect 35866 14260 35894 14368
rect 36081 14365 36093 14368
rect 36127 14365 36139 14399
rect 36081 14359 36139 14365
rect 36262 14260 36268 14272
rect 35584 14232 35894 14260
rect 36223 14232 36268 14260
rect 35584 14220 35590 14232
rect 36262 14220 36268 14232
rect 36320 14220 36326 14272
rect 1104 14170 36892 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 36892 14170
rect 1104 14096 36892 14118
rect 3970 14056 3976 14068
rect 1688 14028 3976 14056
rect 1688 13929 1716 14028
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 5166 14056 5172 14068
rect 4908 14028 5172 14056
rect 1854 13948 1860 14000
rect 1912 13988 1918 14000
rect 1949 13991 2007 13997
rect 1949 13988 1961 13991
rect 1912 13960 1961 13988
rect 1912 13948 1918 13960
rect 1949 13957 1961 13960
rect 1995 13957 2007 13991
rect 4908 13988 4936 14028
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 11057 14059 11115 14065
rect 6880 14028 10548 14056
rect 6880 14016 6886 14028
rect 7006 13988 7012 14000
rect 3174 13960 4936 13988
rect 5750 13960 7012 13988
rect 1949 13951 2007 13957
rect 7006 13948 7012 13960
rect 7064 13948 7070 14000
rect 7374 13988 7380 14000
rect 7335 13960 7380 13988
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 9674 13988 9680 14000
rect 8602 13960 9680 13988
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 9766 13948 9772 14000
rect 9824 13988 9830 14000
rect 9861 13991 9919 13997
rect 9861 13988 9873 13991
rect 9824 13960 9873 13988
rect 9824 13948 9830 13960
rect 9861 13957 9873 13960
rect 9907 13957 9919 13991
rect 9861 13951 9919 13957
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 4028 13892 4261 13920
rect 4028 13880 4034 13892
rect 4249 13889 4261 13892
rect 4295 13889 4307 13923
rect 9950 13920 9956 13932
rect 4249 13883 4307 13889
rect 5736 13892 6868 13920
rect 2038 13812 2044 13864
rect 2096 13852 2102 13864
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 2096 13824 3433 13852
rect 2096 13812 2102 13824
rect 3421 13821 3433 13824
rect 3467 13821 3479 13855
rect 4522 13852 4528 13864
rect 4483 13824 4528 13852
rect 3421 13815 3479 13821
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 4614 13812 4620 13864
rect 4672 13852 4678 13864
rect 5736 13852 5764 13892
rect 5994 13852 6000 13864
rect 4672 13824 5764 13852
rect 5955 13824 6000 13852
rect 4672 13812 4678 13824
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 6638 13784 6644 13796
rect 6599 13756 6644 13784
rect 6638 13744 6644 13756
rect 6696 13744 6702 13796
rect 6840 13784 6868 13892
rect 8588 13892 9260 13920
rect 9863 13892 9956 13920
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 6972 13824 7113 13852
rect 6972 13812 6978 13824
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 8588 13852 8616 13892
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 7101 13815 7159 13821
rect 7208 13824 8616 13852
rect 8680 13824 9137 13852
rect 7208 13784 7236 13824
rect 6840 13756 7236 13784
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 8680 13716 8708 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 9232 13852 9260 13892
rect 9950 13880 9956 13892
rect 10008 13920 10014 13932
rect 10410 13920 10416 13932
rect 10008 13892 10416 13920
rect 10008 13880 10014 13892
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 10520 13920 10548 14028
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 11974 14056 11980 14068
rect 11103 14028 11980 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12069 14059 12127 14065
rect 12069 14025 12081 14059
rect 12115 14056 12127 14059
rect 14366 14056 14372 14068
rect 12115 14028 14372 14056
rect 12115 14025 12127 14028
rect 12069 14019 12127 14025
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 21085 14059 21143 14065
rect 21085 14025 21097 14059
rect 21131 14056 21143 14059
rect 22462 14056 22468 14068
rect 21131 14028 22468 14056
rect 21131 14025 21143 14028
rect 21085 14019 21143 14025
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 12802 13988 12808 14000
rect 12763 13960 12808 13988
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 14274 13988 14280 14000
rect 14235 13960 14280 13988
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14826 13988 14832 14000
rect 14787 13960 14832 13988
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 15470 13988 15476 14000
rect 15431 13960 15476 13988
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 15562 13948 15568 14000
rect 15620 13988 15626 14000
rect 16945 13991 17003 13997
rect 16945 13988 16957 13991
rect 15620 13960 16957 13988
rect 15620 13948 15626 13960
rect 16945 13957 16957 13960
rect 16991 13957 17003 13991
rect 16945 13951 17003 13957
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 18509 13991 18567 13997
rect 18509 13988 18521 13991
rect 17083 13960 18521 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 18509 13957 18521 13960
rect 18555 13957 18567 13991
rect 19978 13988 19984 14000
rect 18509 13951 18567 13957
rect 18616 13960 19984 13988
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10520 13892 10977 13920
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 11992 13852 12020 13883
rect 17678 13880 17684 13932
rect 17736 13920 17742 13932
rect 17862 13920 17868 13932
rect 17736 13892 17868 13920
rect 17736 13880 17742 13892
rect 17862 13880 17868 13892
rect 17920 13880 17926 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18616 13929 18644 13960
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 20349 13991 20407 13997
rect 20349 13957 20361 13991
rect 20395 13988 20407 13991
rect 22094 13988 22100 14000
rect 20395 13960 21312 13988
rect 22055 13960 22100 13988
rect 20395 13957 20407 13960
rect 20349 13951 20407 13957
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18472 13892 18613 13920
rect 18472 13880 18478 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 18782 13880 18788 13932
rect 18840 13920 18846 13932
rect 19245 13923 19303 13929
rect 19245 13920 19257 13923
rect 18840 13892 19257 13920
rect 18840 13880 18846 13892
rect 19245 13889 19257 13892
rect 19291 13889 19303 13923
rect 20990 13920 20996 13932
rect 20951 13892 20996 13920
rect 19245 13883 19303 13889
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 9232 13824 12020 13852
rect 9125 13815 9183 13821
rect 9140 13784 9168 13815
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 12308 13824 12725 13852
rect 12308 13812 12314 13824
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 13354 13852 13360 13864
rect 13315 13824 13360 13852
rect 12713 13815 12771 13821
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 14182 13852 14188 13864
rect 14143 13824 14188 13852
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 15102 13812 15108 13864
rect 15160 13852 15166 13864
rect 15381 13855 15439 13861
rect 15381 13852 15393 13855
rect 15160 13824 15393 13852
rect 15160 13812 15166 13824
rect 15381 13821 15393 13824
rect 15427 13821 15439 13855
rect 15381 13815 15439 13821
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13852 16083 13855
rect 17402 13852 17408 13864
rect 16071 13824 17408 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13852 17647 13855
rect 19797 13855 19855 13861
rect 19797 13852 19809 13855
rect 17635 13824 19809 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 19260 13796 19288 13824
rect 19797 13821 19809 13824
rect 19843 13821 19855 13855
rect 19797 13815 19855 13821
rect 20162 13812 20168 13864
rect 20220 13852 20226 13864
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 20220 13824 20453 13852
rect 20220 13812 20226 13824
rect 20441 13821 20453 13824
rect 20487 13821 20499 13855
rect 21284 13852 21312 13960
rect 22094 13948 22100 13960
rect 22152 13948 22158 14000
rect 22189 13991 22247 13997
rect 22189 13957 22201 13991
rect 22235 13988 22247 13991
rect 23293 13991 23351 13997
rect 23293 13988 23305 13991
rect 22235 13960 23305 13988
rect 22235 13957 22247 13960
rect 22189 13951 22247 13957
rect 23293 13957 23305 13960
rect 23339 13957 23351 13991
rect 23293 13951 23351 13957
rect 23474 13948 23480 14000
rect 23532 13988 23538 14000
rect 32398 13988 32404 14000
rect 23532 13960 32404 13988
rect 23532 13948 23538 13960
rect 32398 13948 32404 13960
rect 32456 13948 32462 14000
rect 22738 13880 22744 13932
rect 22796 13920 22802 13932
rect 23382 13920 23388 13932
rect 22796 13892 22841 13920
rect 23343 13892 23388 13920
rect 22796 13880 22802 13892
rect 23382 13880 23388 13892
rect 23440 13920 23446 13932
rect 23845 13923 23903 13929
rect 23845 13920 23857 13923
rect 23440 13892 23857 13920
rect 23440 13880 23446 13892
rect 23845 13889 23857 13892
rect 23891 13889 23903 13923
rect 23845 13883 23903 13889
rect 22462 13852 22468 13864
rect 21284 13824 22468 13852
rect 20441 13815 20499 13821
rect 22462 13812 22468 13824
rect 22520 13812 22526 13864
rect 9398 13784 9404 13796
rect 9140 13756 9404 13784
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 9490 13744 9496 13796
rect 9548 13784 9554 13796
rect 12894 13784 12900 13796
rect 9548 13756 12900 13784
rect 9548 13744 9554 13756
rect 12894 13744 12900 13756
rect 12952 13744 12958 13796
rect 19242 13744 19248 13796
rect 19300 13744 19306 13796
rect 3568 13688 8708 13716
rect 10505 13719 10563 13725
rect 3568 13676 3574 13688
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 10594 13716 10600 13728
rect 10551 13688 10600 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 18966 13716 18972 13728
rect 11204 13688 18972 13716
rect 11204 13676 11210 13688
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 19150 13716 19156 13728
rect 19111 13688 19156 13716
rect 19150 13676 19156 13688
rect 19208 13676 19214 13728
rect 1104 13626 36892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 36892 13626
rect 1104 13552 36892 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 1946 13512 1952 13524
rect 1719 13484 1952 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 1946 13472 1952 13484
rect 2004 13512 2010 13524
rect 2406 13512 2412 13524
rect 2004 13484 2412 13512
rect 2004 13472 2010 13484
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 4982 13512 4988 13524
rect 4764 13484 4988 13512
rect 4764 13472 4770 13484
rect 4982 13472 4988 13484
rect 5040 13512 5046 13524
rect 5040 13484 5764 13512
rect 5040 13472 5046 13484
rect 4798 13404 4804 13456
rect 4856 13444 4862 13456
rect 5442 13444 5448 13456
rect 4856 13416 5448 13444
rect 4856 13404 4862 13416
rect 5442 13404 5448 13416
rect 5500 13404 5506 13456
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13413 5687 13447
rect 5736 13444 5764 13484
rect 6638 13472 6644 13524
rect 6696 13512 6702 13524
rect 8846 13512 8852 13524
rect 6696 13484 8852 13512
rect 6696 13472 6702 13484
rect 8846 13472 8852 13484
rect 8904 13512 8910 13524
rect 9122 13512 9128 13524
rect 8904 13484 9128 13512
rect 8904 13472 8910 13484
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 9769 13515 9827 13521
rect 9769 13512 9781 13515
rect 9272 13484 9781 13512
rect 9272 13472 9278 13484
rect 9769 13481 9781 13484
rect 9815 13481 9827 13515
rect 9769 13475 9827 13481
rect 13633 13515 13691 13521
rect 13633 13481 13645 13515
rect 13679 13512 13691 13515
rect 14274 13512 14280 13524
rect 13679 13484 14280 13512
rect 13679 13481 13691 13484
rect 13633 13475 13691 13481
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 15197 13515 15255 13521
rect 15197 13481 15209 13515
rect 15243 13512 15255 13515
rect 15378 13512 15384 13524
rect 15243 13484 15384 13512
rect 15243 13481 15255 13484
rect 15197 13475 15255 13481
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 16209 13515 16267 13521
rect 16209 13512 16221 13515
rect 15528 13484 16221 13512
rect 15528 13472 15534 13484
rect 16209 13481 16221 13484
rect 16255 13481 16267 13515
rect 16209 13475 16267 13481
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18049 13515 18107 13521
rect 18049 13512 18061 13515
rect 18012 13484 18061 13512
rect 18012 13472 18018 13484
rect 18049 13481 18061 13484
rect 18095 13481 18107 13515
rect 18049 13475 18107 13481
rect 18782 13472 18788 13524
rect 18840 13512 18846 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 18840 13484 19441 13512
rect 18840 13472 18846 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 20070 13472 20076 13524
rect 20128 13512 20134 13524
rect 20165 13515 20223 13521
rect 20165 13512 20177 13515
rect 20128 13484 20177 13512
rect 20128 13472 20134 13484
rect 20165 13481 20177 13484
rect 20211 13481 20223 13515
rect 20165 13475 20223 13481
rect 21634 13472 21640 13524
rect 21692 13512 21698 13524
rect 21821 13515 21879 13521
rect 21821 13512 21833 13515
rect 21692 13484 21833 13512
rect 21692 13472 21698 13484
rect 21821 13481 21833 13484
rect 21867 13481 21879 13515
rect 22462 13512 22468 13524
rect 22423 13484 22468 13512
rect 21821 13475 21879 13481
rect 22462 13472 22468 13484
rect 22520 13472 22526 13524
rect 5736 13416 6684 13444
rect 5629 13407 5687 13413
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13376 3479 13379
rect 5644 13376 5672 13407
rect 6454 13376 6460 13388
rect 3467 13348 6460 13376
rect 3467 13345 3479 13348
rect 3421 13339 3479 13345
rect 6454 13336 6460 13348
rect 6512 13376 6518 13388
rect 6549 13379 6607 13385
rect 6549 13376 6561 13379
rect 6512 13348 6561 13376
rect 6512 13336 6518 13348
rect 6549 13345 6561 13348
rect 6595 13345 6607 13379
rect 6656 13376 6684 13416
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 8168 13416 10425 13444
rect 8168 13404 8174 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 10413 13407 10471 13413
rect 13538 13404 13544 13456
rect 13596 13404 13602 13456
rect 14553 13447 14611 13453
rect 14553 13413 14565 13447
rect 14599 13444 14611 13447
rect 15286 13444 15292 13456
rect 14599 13416 15292 13444
rect 14599 13413 14611 13416
rect 14553 13407 14611 13413
rect 15286 13404 15292 13416
rect 15344 13404 15350 13456
rect 18966 13404 18972 13456
rect 19024 13444 19030 13456
rect 20806 13444 20812 13456
rect 19024 13416 20812 13444
rect 19024 13404 19030 13416
rect 20806 13404 20812 13416
rect 20864 13444 20870 13456
rect 20990 13444 20996 13456
rect 20864 13416 20996 13444
rect 20864 13404 20870 13416
rect 20990 13404 20996 13416
rect 21048 13404 21054 13456
rect 8573 13379 8631 13385
rect 6656 13348 8064 13376
rect 6549 13339 6607 13345
rect 4341 13311 4399 13317
rect 4341 13277 4353 13311
rect 4387 13308 4399 13311
rect 5350 13308 5356 13320
rect 4387 13280 5356 13308
rect 4387 13277 4399 13280
rect 4341 13271 4399 13277
rect 5350 13268 5356 13280
rect 5408 13308 5414 13320
rect 5534 13308 5540 13320
rect 5408 13280 5540 13308
rect 5408 13268 5414 13280
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 8036 13308 8064 13348
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 8662 13376 8668 13388
rect 8619 13348 8668 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 11146 13376 11152 13388
rect 8772 13348 11152 13376
rect 8772 13308 8800 13348
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 13556 13376 13584 13404
rect 16758 13376 16764 13388
rect 13556 13348 15148 13376
rect 5684 13280 6592 13308
rect 8036 13280 8800 13308
rect 9861 13311 9919 13317
rect 5684 13268 5690 13280
rect 3145 13243 3203 13249
rect 2714 13212 2774 13240
rect 2746 13172 2774 13212
rect 3145 13209 3157 13243
rect 3191 13240 3203 13243
rect 5994 13240 6000 13252
rect 3191 13212 6000 13240
rect 3191 13209 3203 13212
rect 3145 13203 3203 13209
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 6564 13240 6592 13280
rect 9861 13277 9873 13311
rect 9907 13308 9919 13311
rect 9950 13308 9956 13320
rect 9907 13280 9956 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 10468 13280 10517 13308
rect 10468 13268 10474 13280
rect 10505 13277 10517 13280
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11425 13311 11483 13317
rect 11425 13308 11437 13311
rect 11388 13280 11437 13308
rect 11388 13268 11394 13280
rect 11425 13277 11437 13280
rect 11471 13308 11483 13311
rect 11514 13308 11520 13320
rect 11471 13280 11520 13308
rect 11471 13277 11483 13280
rect 11425 13271 11483 13277
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 13541 13311 13599 13317
rect 13541 13308 13553 13311
rect 13504 13280 13553 13308
rect 13504 13268 13510 13280
rect 13541 13277 13553 13280
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 15120 13317 15148 13348
rect 16316 13348 16764 13376
rect 16316 13317 16344 13348
rect 16758 13336 16764 13348
rect 16816 13376 16822 13388
rect 20898 13376 20904 13388
rect 16816 13348 18000 13376
rect 16816 13336 16822 13348
rect 17972 13317 18000 13348
rect 18800 13348 20904 13376
rect 18800 13320 18828 13348
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 13872 13280 14473 13308
rect 13872 13268 13878 13280
rect 14461 13277 14473 13280
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 16301 13311 16359 13317
rect 16301 13277 16313 13311
rect 16347 13277 16359 13311
rect 16301 13271 16359 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13277 18015 13311
rect 18782 13308 18788 13320
rect 18743 13280 18788 13308
rect 17957 13271 18015 13277
rect 18782 13268 18788 13280
rect 18840 13268 18846 13320
rect 19978 13268 19984 13320
rect 20036 13308 20042 13320
rect 20073 13311 20131 13317
rect 20073 13308 20085 13311
rect 20036 13280 20085 13308
rect 20036 13268 20042 13280
rect 20073 13277 20085 13280
rect 20119 13277 20131 13311
rect 20073 13271 20131 13277
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13308 21971 13311
rect 22186 13308 22192 13320
rect 21959 13280 22192 13308
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 22186 13268 22192 13280
rect 22244 13308 22250 13320
rect 22557 13311 22615 13317
rect 22557 13308 22569 13311
rect 22244 13280 22569 13308
rect 22244 13268 22250 13280
rect 22557 13277 22569 13280
rect 22603 13308 22615 13311
rect 23017 13311 23075 13317
rect 23017 13308 23029 13311
rect 22603 13280 23029 13308
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 23017 13277 23029 13280
rect 23063 13308 23075 13311
rect 23382 13308 23388 13320
rect 23063 13280 23388 13308
rect 23063 13277 23075 13280
rect 23017 13271 23075 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 35894 13268 35900 13320
rect 35952 13308 35958 13320
rect 35952 13280 35997 13308
rect 35952 13268 35958 13280
rect 6564 13212 6776 13240
rect 6454 13172 6460 13184
rect 2746 13144 6460 13172
rect 6454 13132 6460 13144
rect 6512 13132 6518 13184
rect 6748 13172 6776 13212
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 6880 13212 6925 13240
rect 6880 13200 6886 13212
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 9122 13240 9128 13252
rect 7156 13212 7314 13240
rect 9083 13212 9128 13240
rect 7156 13200 7162 13212
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 12158 13240 12164 13252
rect 12119 13212 12164 13240
rect 12158 13200 12164 13212
rect 12216 13200 12222 13252
rect 12253 13243 12311 13249
rect 12253 13209 12265 13243
rect 12299 13209 12311 13243
rect 12253 13203 12311 13209
rect 12805 13243 12863 13249
rect 12805 13209 12817 13243
rect 12851 13240 12863 13243
rect 13170 13240 13176 13252
rect 12851 13212 13176 13240
rect 12851 13209 12863 13212
rect 12805 13203 12863 13209
rect 9950 13172 9956 13184
rect 6748 13144 9956 13172
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 11517 13175 11575 13181
rect 11517 13141 11529 13175
rect 11563 13172 11575 13175
rect 12268 13172 12296 13203
rect 13170 13200 13176 13212
rect 13228 13240 13234 13252
rect 13722 13240 13728 13252
rect 13228 13212 13728 13240
rect 13228 13200 13234 13212
rect 13722 13200 13728 13212
rect 13780 13200 13786 13252
rect 11563 13144 12296 13172
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 12342 13132 12348 13184
rect 12400 13172 12406 13184
rect 13832 13172 13860 13268
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 16761 13243 16819 13249
rect 16761 13240 16773 13243
rect 14976 13212 16773 13240
rect 14976 13200 14982 13212
rect 16761 13209 16773 13212
rect 16807 13240 16819 13243
rect 17218 13240 17224 13252
rect 16807 13212 17224 13240
rect 16807 13209 16819 13212
rect 16761 13203 16819 13209
rect 17218 13200 17224 13212
rect 17276 13200 17282 13252
rect 17313 13243 17371 13249
rect 17313 13209 17325 13243
rect 17359 13209 17371 13243
rect 17313 13203 17371 13209
rect 12400 13144 13860 13172
rect 17328 13172 17356 13203
rect 17402 13200 17408 13252
rect 17460 13240 17466 13252
rect 18693 13243 18751 13249
rect 17460 13212 17505 13240
rect 17460 13200 17466 13212
rect 18693 13209 18705 13243
rect 18739 13209 18751 13243
rect 18693 13203 18751 13209
rect 18708 13172 18736 13203
rect 36078 13172 36084 13184
rect 17328 13144 18736 13172
rect 36039 13144 36084 13172
rect 12400 13132 12406 13144
rect 36078 13132 36084 13144
rect 36136 13132 36142 13184
rect 1104 13082 36892 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 36892 13082
rect 1104 13008 36892 13030
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 5813 12971 5871 12977
rect 3016 12940 5672 12968
rect 3016 12928 3022 12940
rect 2866 12860 2872 12912
rect 2924 12860 2930 12912
rect 4341 12903 4399 12909
rect 4341 12869 4353 12903
rect 4387 12900 4399 12903
rect 4614 12900 4620 12912
rect 4387 12872 4620 12900
rect 4387 12869 4399 12872
rect 4341 12863 4399 12869
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 5644 12900 5672 12940
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 7742 12968 7748 12980
rect 5859 12940 7748 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 7926 12928 7932 12980
rect 7984 12968 7990 12980
rect 9490 12968 9496 12980
rect 7984 12940 8892 12968
rect 7984 12928 7990 12940
rect 5644 12872 8050 12900
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12832 3663 12835
rect 3970 12832 3976 12844
rect 3651 12804 3976 12832
rect 3651 12801 3663 12804
rect 3605 12795 3663 12801
rect 3970 12792 3976 12804
rect 4028 12832 4034 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 4028 12804 4077 12832
rect 4028 12792 4034 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 5442 12792 5448 12844
rect 5500 12792 5506 12844
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6788 12804 6837 12832
rect 6788 12792 6794 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 8864 12832 8892 12940
rect 9324 12940 9496 12968
rect 9324 12909 9352 12940
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 9950 12968 9956 12980
rect 9911 12940 9956 12968
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10560 12940 10609 12968
rect 10560 12928 10566 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 12437 12971 12495 12977
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 12802 12968 12808 12980
rect 12483 12940 12808 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 12894 12928 12900 12980
rect 12952 12968 12958 12980
rect 12952 12940 15608 12968
rect 12952 12928 12958 12940
rect 9309 12903 9367 12909
rect 9309 12869 9321 12903
rect 9355 12869 9367 12903
rect 9309 12863 9367 12869
rect 9398 12860 9404 12912
rect 9456 12900 9462 12912
rect 13170 12900 13176 12912
rect 9456 12872 12388 12900
rect 13131 12872 13176 12900
rect 9456 12860 9462 12872
rect 9950 12832 9956 12844
rect 8864 12804 9956 12832
rect 6825 12795 6883 12801
rect 9950 12792 9956 12804
rect 10008 12832 10014 12844
rect 12360 12841 12388 12872
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 14366 12900 14372 12912
rect 14327 12872 14372 12900
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 10008 12804 10057 12832
rect 10008 12792 10014 12804
rect 10045 12801 10057 12804
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 12345 12835 12403 12841
rect 12345 12801 12357 12835
rect 12391 12801 12403 12835
rect 12345 12795 12403 12801
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12764 1639 12767
rect 2314 12764 2320 12776
rect 1627 12736 2320 12764
rect 1627 12733 1639 12736
rect 1581 12727 1639 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 3329 12767 3387 12773
rect 3329 12733 3341 12767
rect 3375 12764 3387 12767
rect 3694 12764 3700 12776
rect 3375 12736 3700 12764
rect 3375 12733 3387 12736
rect 3329 12727 3387 12733
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 4706 12764 4712 12776
rect 3804 12736 4712 12764
rect 2332 12628 2360 12724
rect 3804 12696 3832 12736
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 7282 12764 7288 12776
rect 7243 12736 7288 12764
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 8202 12764 8208 12776
rect 7607 12736 8208 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 10520 12764 10548 12795
rect 9548 12736 10548 12764
rect 9548 12724 9554 12736
rect 3528 12668 3832 12696
rect 3528 12628 3556 12668
rect 5718 12656 5724 12708
rect 5776 12696 5782 12708
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 5776 12668 6653 12696
rect 5776 12656 5782 12668
rect 6641 12665 6653 12668
rect 6687 12665 6699 12699
rect 6641 12659 6699 12665
rect 8662 12656 8668 12708
rect 8720 12696 8726 12708
rect 11716 12696 11744 12795
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12764 13139 12767
rect 13998 12764 14004 12776
rect 13127 12736 14004 12764
rect 13127 12733 13139 12736
rect 13081 12727 13139 12733
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14274 12764 14280 12776
rect 14235 12736 14280 12764
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14553 12767 14611 12773
rect 14553 12733 14565 12767
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 8720 12668 11744 12696
rect 11793 12699 11851 12705
rect 8720 12656 8726 12668
rect 11793 12665 11805 12699
rect 11839 12696 11851 12699
rect 12986 12696 12992 12708
rect 11839 12668 12992 12696
rect 11839 12665 11851 12668
rect 11793 12659 11851 12665
rect 12986 12656 12992 12668
rect 13044 12656 13050 12708
rect 13354 12656 13360 12708
rect 13412 12696 13418 12708
rect 13633 12699 13691 12705
rect 13633 12696 13645 12699
rect 13412 12668 13645 12696
rect 13412 12656 13418 12668
rect 13633 12665 13645 12668
rect 13679 12665 13691 12699
rect 13633 12659 13691 12665
rect 2332 12600 3556 12628
rect 3602 12588 3608 12640
rect 3660 12628 3666 12640
rect 6546 12628 6552 12640
rect 3660 12600 6552 12628
rect 3660 12588 3666 12600
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 13648 12628 13676 12659
rect 13722 12656 13728 12708
rect 13780 12696 13786 12708
rect 14568 12696 14596 12727
rect 13780 12668 14596 12696
rect 13780 12656 13786 12668
rect 15378 12628 15384 12640
rect 13648 12600 15384 12628
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 15580 12628 15608 12940
rect 17402 12928 17408 12980
rect 17460 12968 17466 12980
rect 20809 12971 20867 12977
rect 20809 12968 20821 12971
rect 17460 12940 20821 12968
rect 17460 12928 17466 12940
rect 20809 12937 20821 12940
rect 20855 12937 20867 12971
rect 20809 12931 20867 12937
rect 22097 12971 22155 12977
rect 22097 12937 22109 12971
rect 22143 12968 22155 12971
rect 22186 12968 22192 12980
rect 22143 12940 22192 12968
rect 22143 12937 22155 12940
rect 22097 12931 22155 12937
rect 22186 12928 22192 12940
rect 22244 12928 22250 12980
rect 16117 12903 16175 12909
rect 16117 12869 16129 12903
rect 16163 12900 16175 12903
rect 16666 12900 16672 12912
rect 16163 12872 16672 12900
rect 16163 12869 16175 12872
rect 16117 12863 16175 12869
rect 16666 12860 16672 12872
rect 16724 12860 16730 12912
rect 17037 12903 17095 12909
rect 17037 12869 17049 12903
rect 17083 12900 17095 12903
rect 19150 12900 19156 12912
rect 17083 12872 19156 12900
rect 17083 12869 17095 12872
rect 17037 12863 17095 12869
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 19426 12900 19432 12912
rect 19387 12872 19432 12900
rect 19426 12860 19432 12872
rect 19484 12860 19490 12912
rect 19521 12903 19579 12909
rect 19521 12869 19533 12903
rect 19567 12900 19579 12903
rect 20254 12900 20260 12912
rect 19567 12872 20260 12900
rect 19567 12869 19579 12872
rect 19521 12863 19579 12869
rect 20254 12860 20260 12872
rect 20312 12900 20318 12912
rect 20530 12900 20536 12912
rect 20312 12872 20536 12900
rect 20312 12860 20318 12872
rect 20530 12860 20536 12872
rect 20588 12860 20594 12912
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12832 18107 12835
rect 18322 12832 18328 12844
rect 18095 12804 18328 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 19978 12792 19984 12844
rect 20036 12832 20042 12844
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 20036 12804 20085 12832
rect 20036 12792 20042 12804
rect 20073 12801 20085 12804
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 20901 12835 20959 12841
rect 20901 12801 20913 12835
rect 20947 12832 20959 12835
rect 35621 12835 35679 12841
rect 20947 12804 21496 12832
rect 20947 12801 20959 12804
rect 20901 12795 20959 12801
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12733 15991 12767
rect 16206 12764 16212 12776
rect 16119 12736 16212 12764
rect 15933 12727 15991 12733
rect 15948 12696 15976 12727
rect 16206 12724 16212 12736
rect 16264 12764 16270 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16264 12736 16957 12764
rect 16264 12724 16270 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 17218 12764 17224 12776
rect 17179 12736 17224 12764
rect 16945 12727 17003 12733
rect 17218 12724 17224 12736
rect 17276 12724 17282 12776
rect 18138 12724 18144 12776
rect 18196 12764 18202 12776
rect 19242 12764 19248 12776
rect 18196 12736 19248 12764
rect 18196 12724 18202 12736
rect 19242 12724 19248 12736
rect 19300 12724 19306 12776
rect 16574 12696 16580 12708
rect 15948 12668 16580 12696
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 21468 12705 21496 12804
rect 35621 12801 35633 12835
rect 35667 12832 35679 12835
rect 35802 12832 35808 12844
rect 35667 12804 35808 12832
rect 35667 12801 35679 12804
rect 35621 12795 35679 12801
rect 35802 12792 35808 12804
rect 35860 12832 35866 12844
rect 36265 12835 36323 12841
rect 36265 12832 36277 12835
rect 35860 12804 36277 12832
rect 35860 12792 35866 12804
rect 36265 12801 36277 12804
rect 36311 12801 36323 12835
rect 36265 12795 36323 12801
rect 21453 12699 21511 12705
rect 21453 12665 21465 12699
rect 21499 12696 21511 12699
rect 22094 12696 22100 12708
rect 21499 12668 22100 12696
rect 21499 12665 21511 12668
rect 21453 12659 21511 12665
rect 22094 12656 22100 12668
rect 22152 12696 22158 12708
rect 36081 12699 36139 12705
rect 36081 12696 36093 12699
rect 22152 12668 36093 12696
rect 22152 12656 22158 12668
rect 36081 12665 36093 12668
rect 36127 12665 36139 12699
rect 36081 12659 36139 12665
rect 18782 12628 18788 12640
rect 15580 12600 18788 12628
rect 18782 12588 18788 12600
rect 18840 12628 18846 12640
rect 18966 12628 18972 12640
rect 18840 12600 18972 12628
rect 18840 12588 18846 12600
rect 18966 12588 18972 12600
rect 19024 12588 19030 12640
rect 20070 12588 20076 12640
rect 20128 12628 20134 12640
rect 20165 12631 20223 12637
rect 20165 12628 20177 12631
rect 20128 12600 20177 12628
rect 20128 12588 20134 12600
rect 20165 12597 20177 12600
rect 20211 12597 20223 12631
rect 20165 12591 20223 12597
rect 1104 12538 36892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 36892 12538
rect 1104 12464 36892 12486
rect 1673 12427 1731 12433
rect 1673 12393 1685 12427
rect 1719 12424 1731 12427
rect 1854 12424 1860 12436
rect 1719 12396 1860 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 1854 12384 1860 12396
rect 1912 12424 1918 12436
rect 2498 12424 2504 12436
rect 1912 12396 2504 12424
rect 1912 12384 1918 12396
rect 2498 12384 2504 12396
rect 2556 12384 2562 12436
rect 5350 12424 5356 12436
rect 4724 12396 5356 12424
rect 4724 12356 4752 12396
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 9306 12424 9312 12436
rect 6052 12396 8524 12424
rect 9267 12396 9312 12424
rect 6052 12384 6058 12396
rect 6730 12356 6736 12368
rect 4356 12328 4752 12356
rect 5920 12328 6736 12356
rect 3145 12291 3203 12297
rect 3145 12257 3157 12291
rect 3191 12288 3203 12291
rect 4356 12288 4384 12328
rect 5920 12288 5948 12328
rect 6730 12316 6736 12328
rect 6788 12316 6794 12368
rect 8496 12356 8524 12396
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 9953 12427 10011 12433
rect 9953 12424 9965 12427
rect 9916 12396 9965 12424
rect 9916 12384 9922 12396
rect 9953 12393 9965 12396
rect 9999 12393 10011 12427
rect 9953 12387 10011 12393
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 10962 12424 10968 12436
rect 10643 12396 10968 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 13630 12424 13636 12436
rect 13591 12396 13636 12424
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 14366 12424 14372 12436
rect 14327 12396 14372 12424
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 15930 12424 15936 12436
rect 15488 12396 15936 12424
rect 8496 12328 10548 12356
rect 3191 12260 4384 12288
rect 4448 12260 5948 12288
rect 5997 12291 6055 12297
rect 3191 12257 3203 12260
rect 3145 12251 3203 12257
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 3970 12220 3976 12232
rect 3467 12192 3976 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 3970 12180 3976 12192
rect 4028 12180 4034 12232
rect 4448 12152 4476 12260
rect 5997 12257 6009 12291
rect 6043 12288 6055 12291
rect 6914 12288 6920 12300
rect 6043 12260 6920 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 8573 12291 8631 12297
rect 8573 12288 8585 12291
rect 7340 12260 8585 12288
rect 7340 12248 7346 12260
rect 8573 12257 8585 12260
rect 8619 12257 8631 12291
rect 8573 12251 8631 12257
rect 8662 12248 8668 12300
rect 8720 12288 8726 12300
rect 9858 12288 9864 12300
rect 8720 12260 9864 12288
rect 8720 12248 8726 12260
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 6822 12220 6828 12232
rect 6420 12192 6828 12220
rect 6420 12180 6426 12192
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 8812 12192 9413 12220
rect 8812 12180 8818 12192
rect 9401 12189 9413 12192
rect 9447 12220 9459 12223
rect 9490 12220 9496 12232
rect 9447 12192 9496 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 9490 12180 9496 12192
rect 9548 12180 9554 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9950 12220 9956 12232
rect 9824 12192 9956 12220
rect 9824 12180 9830 12192
rect 9950 12180 9956 12192
rect 10008 12220 10014 12232
rect 10520 12229 10548 12328
rect 11164 12328 12020 12356
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 10008 12192 10057 12220
rect 10008 12180 10014 12192
rect 10045 12189 10057 12192
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12189 10563 12223
rect 10505 12183 10563 12189
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 11164 12220 11192 12328
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12288 11575 12291
rect 11606 12288 11612 12300
rect 11563 12260 11612 12288
rect 11563 12257 11575 12260
rect 11517 12251 11575 12257
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 11756 12260 11805 12288
rect 11756 12248 11762 12260
rect 11793 12257 11805 12260
rect 11839 12257 11851 12291
rect 11793 12251 11851 12257
rect 10744 12192 11192 12220
rect 10744 12180 10750 12192
rect 2714 12124 4476 12152
rect 5290 12124 5672 12152
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 5350 12084 5356 12096
rect 4295 12056 5356 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5644 12084 5672 12124
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 6549 12155 6607 12161
rect 5776 12124 5821 12152
rect 5776 12112 5782 12124
rect 6549 12121 6561 12155
rect 6595 12152 6607 12155
rect 8297 12155 8355 12161
rect 6595 12124 7052 12152
rect 7866 12124 8248 12152
rect 6595 12121 6607 12124
rect 6549 12115 6607 12121
rect 6914 12084 6920 12096
rect 5644 12056 6920 12084
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 7024 12084 7052 12124
rect 8018 12084 8024 12096
rect 7024 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8220 12084 8248 12124
rect 8297 12121 8309 12155
rect 8343 12152 8355 12155
rect 8386 12152 8392 12164
rect 8343 12124 8392 12152
rect 8343 12121 8355 12124
rect 8297 12115 8355 12121
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 11422 12152 11428 12164
rect 8720 12124 11428 12152
rect 8720 12112 8726 12124
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 11701 12155 11759 12161
rect 11701 12121 11713 12155
rect 11747 12121 11759 12155
rect 11992 12152 12020 12328
rect 13998 12316 14004 12368
rect 14056 12356 14062 12368
rect 15488 12356 15516 12396
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 16666 12424 16672 12436
rect 16627 12396 16672 12424
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 16850 12384 16856 12436
rect 16908 12424 16914 12436
rect 18509 12427 18567 12433
rect 16908 12396 18000 12424
rect 16908 12384 16914 12396
rect 17402 12356 17408 12368
rect 14056 12328 15516 12356
rect 15580 12328 17408 12356
rect 14056 12316 14062 12328
rect 12066 12248 12072 12300
rect 12124 12288 12130 12300
rect 15580 12297 15608 12328
rect 17402 12316 17408 12328
rect 17460 12356 17466 12368
rect 17972 12356 18000 12396
rect 18509 12393 18521 12427
rect 18555 12424 18567 12427
rect 18966 12424 18972 12436
rect 18555 12396 18972 12424
rect 18555 12393 18567 12396
rect 18509 12387 18567 12393
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 17460 12328 17908 12356
rect 17972 12328 22094 12356
rect 17460 12316 17466 12328
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 12124 12260 14933 12288
rect 12124 12248 12130 12260
rect 14921 12257 14933 12260
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12257 15623 12291
rect 15565 12251 15623 12257
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 17880 12297 17908 12328
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 16632 12260 17233 12288
rect 16632 12248 16638 12260
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 17865 12291 17923 12297
rect 17865 12257 17877 12291
rect 17911 12257 17923 12291
rect 22066 12288 22094 12328
rect 35526 12288 35532 12300
rect 22066 12260 35532 12288
rect 17865 12251 17923 12257
rect 35526 12248 35532 12260
rect 35584 12248 35590 12300
rect 14458 12220 14464 12232
rect 13280 12192 14320 12220
rect 14419 12192 14464 12220
rect 12437 12155 12495 12161
rect 12437 12152 12449 12155
rect 11992 12124 12449 12152
rect 11701 12115 11759 12121
rect 12437 12121 12449 12124
rect 12483 12121 12495 12155
rect 12986 12152 12992 12164
rect 12947 12124 12992 12152
rect 12437 12115 12495 12121
rect 9306 12084 9312 12096
rect 8220 12056 9312 12084
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 10962 12044 10968 12096
rect 11020 12084 11026 12096
rect 11716 12084 11744 12115
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 13081 12155 13139 12161
rect 13081 12121 13093 12155
rect 13127 12152 13139 12155
rect 13280 12152 13308 12192
rect 13127 12124 13308 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 11020 12056 11744 12084
rect 11020 12044 11026 12056
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 13998 12084 14004 12096
rect 11848 12056 14004 12084
rect 11848 12044 11854 12056
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 14292 12084 14320 12192
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 16758 12220 16764 12232
rect 16719 12192 16764 12220
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 15470 12152 15476 12164
rect 15431 12124 15476 12152
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 15620 12124 17724 12152
rect 15620 12112 15626 12124
rect 15654 12084 15660 12096
rect 14292 12056 15660 12084
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 17586 12084 17592 12096
rect 15988 12056 17592 12084
rect 15988 12044 15994 12056
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 17696 12084 17724 12124
rect 17770 12112 17776 12164
rect 17828 12161 17834 12164
rect 17828 12152 17838 12161
rect 19521 12155 19579 12161
rect 19521 12152 19533 12155
rect 17828 12124 17873 12152
rect 19306 12124 19533 12152
rect 17828 12115 17838 12124
rect 17828 12112 17834 12115
rect 19306 12084 19334 12124
rect 19521 12121 19533 12124
rect 19567 12121 19579 12155
rect 20070 12152 20076 12164
rect 20031 12124 20076 12152
rect 19521 12115 19579 12121
rect 17696 12056 19334 12084
rect 19536 12084 19564 12115
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 20165 12155 20223 12161
rect 20165 12121 20177 12155
rect 20211 12152 20223 12155
rect 20717 12155 20775 12161
rect 20717 12152 20729 12155
rect 20211 12124 20729 12152
rect 20211 12121 20223 12124
rect 20165 12115 20223 12121
rect 20717 12121 20729 12124
rect 20763 12121 20775 12155
rect 20717 12115 20775 12121
rect 21082 12084 21088 12096
rect 19536 12056 21088 12084
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 1104 11994 36892 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 36892 11994
rect 1104 11920 36892 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 1670 11880 1676 11892
rect 1627 11852 1676 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 6733 11883 6791 11889
rect 1820 11852 3464 11880
rect 1820 11840 1826 11852
rect 3326 11812 3332 11824
rect 2622 11784 3332 11812
rect 3326 11772 3332 11784
rect 3384 11772 3390 11824
rect 3436 11744 3464 11852
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 7558 11880 7564 11892
rect 6779 11852 7564 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 10042 11880 10048 11892
rect 7668 11852 9076 11880
rect 10003 11852 10048 11880
rect 7668 11812 7696 11852
rect 3804 11784 4738 11812
rect 5552 11784 7696 11812
rect 7745 11815 7803 11821
rect 3804 11744 3832 11784
rect 3436 11716 3832 11744
rect 3053 11679 3111 11685
rect 3053 11645 3065 11679
rect 3099 11676 3111 11679
rect 3329 11679 3387 11685
rect 3099 11648 3280 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 3252 11608 3280 11648
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 3878 11676 3884 11688
rect 3375 11648 3884 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 4249 11679 4307 11685
rect 4249 11645 4261 11679
rect 4295 11676 4307 11679
rect 4706 11676 4712 11688
rect 4295 11648 4712 11676
rect 4295 11645 4307 11648
rect 4249 11639 4307 11645
rect 3510 11608 3516 11620
rect 3252 11580 3516 11608
rect 3510 11568 3516 11580
rect 3568 11568 3574 11620
rect 1670 11500 1676 11552
rect 1728 11540 1734 11552
rect 3988 11540 4016 11639
rect 4706 11636 4712 11648
rect 4764 11676 4770 11688
rect 4982 11676 4988 11688
rect 4764 11648 4988 11676
rect 4764 11636 4770 11648
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 5350 11568 5356 11620
rect 5408 11608 5414 11620
rect 5552 11608 5580 11784
rect 7745 11781 7757 11815
rect 7791 11812 7803 11815
rect 7834 11812 7840 11824
rect 7791 11784 7840 11812
rect 7791 11781 7803 11784
rect 7745 11775 7803 11781
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 8294 11772 8300 11824
rect 8352 11772 8358 11824
rect 9048 11812 9076 11852
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 12713 11883 12771 11889
rect 10152 11852 12434 11880
rect 10152 11812 10180 11852
rect 9048 11784 10180 11812
rect 10318 11772 10324 11824
rect 10376 11812 10382 11824
rect 10870 11812 10876 11824
rect 10376 11784 10876 11812
rect 10376 11772 10382 11784
rect 10870 11772 10876 11784
rect 10928 11772 10934 11824
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 12406 11812 12434 11852
rect 12713 11849 12725 11883
rect 12759 11880 12771 11883
rect 13170 11880 13176 11892
rect 12759 11852 13176 11880
rect 12759 11849 12771 11852
rect 12713 11843 12771 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 14921 11883 14979 11889
rect 14921 11849 14933 11883
rect 14967 11880 14979 11883
rect 15470 11880 15476 11892
rect 14967 11852 15476 11880
rect 14967 11849 14979 11852
rect 14921 11843 14979 11849
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15565 11883 15623 11889
rect 15565 11849 15577 11883
rect 15611 11880 15623 11883
rect 16206 11880 16212 11892
rect 15611 11852 16212 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 17052 11852 18276 11880
rect 17052 11812 17080 11852
rect 11480 11784 11836 11812
rect 12406 11784 13308 11812
rect 11480 11772 11486 11784
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 6328 11716 6653 11744
rect 6328 11704 6334 11716
rect 6641 11713 6653 11716
rect 6687 11744 6699 11747
rect 6822 11744 6828 11756
rect 6687 11716 6828 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 10226 11744 10232 11756
rect 10187 11716 10232 11744
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11744 11207 11747
rect 11698 11744 11704 11756
rect 11195 11716 11704 11744
rect 11195 11713 11207 11716
rect 11149 11707 11207 11713
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 11808 11744 11836 11784
rect 13280 11753 13308 11784
rect 16224 11784 17080 11812
rect 12621 11747 12679 11753
rect 12621 11744 12633 11747
rect 11808 11716 12633 11744
rect 12621 11713 12633 11716
rect 12667 11713 12679 11747
rect 12621 11707 12679 11713
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11713 13323 11747
rect 13265 11707 13323 11713
rect 13998 11704 14004 11756
rect 14056 11744 14062 11756
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 14056 11716 14197 11744
rect 14056 11704 14062 11716
rect 14185 11713 14197 11716
rect 14231 11744 14243 11747
rect 14458 11744 14464 11756
rect 14231 11716 14464 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 14550 11704 14556 11756
rect 14608 11744 14614 11756
rect 14829 11747 14887 11753
rect 14829 11744 14841 11747
rect 14608 11716 14841 11744
rect 14608 11704 14614 11716
rect 14829 11713 14841 11716
rect 14875 11744 14887 11747
rect 15194 11744 15200 11756
rect 14875 11716 15200 11744
rect 14875 11713 14887 11716
rect 14829 11707 14887 11713
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 15470 11744 15476 11756
rect 15431 11716 15476 11744
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 16224 11753 16252 11784
rect 17126 11772 17132 11824
rect 17184 11812 17190 11824
rect 17313 11815 17371 11821
rect 17313 11812 17325 11815
rect 17184 11784 17325 11812
rect 17184 11772 17190 11784
rect 17313 11781 17325 11784
rect 17359 11781 17371 11815
rect 17313 11775 17371 11781
rect 17402 11772 17408 11824
rect 17460 11812 17466 11824
rect 17460 11784 17505 11812
rect 17460 11772 17466 11784
rect 17586 11772 17592 11824
rect 17644 11812 17650 11824
rect 18248 11812 18276 11852
rect 19426 11840 19432 11892
rect 19484 11880 19490 11892
rect 19705 11883 19763 11889
rect 19705 11880 19717 11883
rect 19484 11852 19717 11880
rect 19484 11840 19490 11852
rect 19705 11849 19717 11852
rect 19751 11849 19763 11883
rect 19705 11843 19763 11849
rect 20349 11883 20407 11889
rect 20349 11849 20361 11883
rect 20395 11880 20407 11883
rect 20806 11880 20812 11892
rect 20395 11852 20812 11880
rect 20395 11849 20407 11852
rect 20349 11843 20407 11849
rect 20254 11812 20260 11824
rect 17644 11784 18000 11812
rect 18248 11784 20260 11812
rect 17644 11772 17650 11784
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16482 11744 16488 11756
rect 16347 11716 16488 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 17972 11744 18000 11784
rect 20254 11772 20260 11784
rect 20312 11772 20318 11824
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17972 11716 18613 11744
rect 18601 11713 18613 11716
rect 18647 11744 18659 11747
rect 19061 11747 19119 11753
rect 19061 11744 19073 11747
rect 18647 11716 19073 11744
rect 18647 11713 18659 11716
rect 18601 11707 18659 11713
rect 19061 11713 19073 11716
rect 19107 11713 19119 11747
rect 19061 11707 19119 11713
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11744 19855 11747
rect 20364 11744 20392 11843
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 19843 11716 20392 11744
rect 19843 11713 19855 11716
rect 19797 11707 19855 11713
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11676 6055 11679
rect 6178 11676 6184 11688
rect 6043 11648 6184 11676
rect 6043 11645 6055 11648
rect 5997 11639 6055 11645
rect 6178 11636 6184 11648
rect 6236 11636 6242 11688
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7340 11648 7481 11676
rect 7340 11636 7346 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 9493 11679 9551 11685
rect 9493 11676 9505 11679
rect 7469 11639 7527 11645
rect 7576 11648 9505 11676
rect 5408 11580 5580 11608
rect 5408 11568 5414 11580
rect 5902 11568 5908 11620
rect 5960 11608 5966 11620
rect 7576 11608 7604 11648
rect 9493 11645 9505 11648
rect 9539 11676 9551 11679
rect 11790 11676 11796 11688
rect 9539 11648 11796 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 5960 11580 7604 11608
rect 5960 11568 5966 11580
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 11900 11608 11928 11639
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 16758 11676 16764 11688
rect 12584 11648 16764 11676
rect 12584 11636 12590 11648
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 17586 11636 17592 11688
rect 17644 11676 17650 11688
rect 18230 11676 18236 11688
rect 17644 11648 18236 11676
rect 17644 11636 17650 11648
rect 18230 11636 18236 11648
rect 18288 11636 18294 11688
rect 9272 11580 11928 11608
rect 13357 11611 13415 11617
rect 9272 11568 9278 11580
rect 13357 11577 13369 11611
rect 13403 11608 13415 11611
rect 13403 11580 17816 11608
rect 13403 11577 13415 11580
rect 13357 11571 13415 11577
rect 1728 11512 4016 11540
rect 1728 11500 1734 11512
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 10778 11540 10784 11552
rect 6328 11512 10784 11540
rect 6328 11500 6334 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 14277 11543 14335 11549
rect 14277 11509 14289 11543
rect 14323 11540 14335 11543
rect 14458 11540 14464 11552
rect 14323 11512 14464 11540
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 16850 11540 16856 11552
rect 14608 11512 16856 11540
rect 14608 11500 14614 11512
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17788 11540 17816 11580
rect 17862 11568 17868 11620
rect 17920 11608 17926 11620
rect 17920 11580 17965 11608
rect 17920 11568 17926 11580
rect 18046 11540 18052 11552
rect 17788 11512 18052 11540
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18506 11540 18512 11552
rect 18467 11512 18512 11540
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 1104 11450 36892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 36892 11450
rect 1104 11376 36892 11398
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11336 3479 11339
rect 3602 11336 3608 11348
rect 3467 11308 3608 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 5166 11336 5172 11348
rect 4295 11308 5172 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 5776 11308 10885 11336
rect 5776 11296 5782 11308
rect 10873 11305 10885 11308
rect 10919 11336 10931 11339
rect 12710 11336 12716 11348
rect 10919 11308 12434 11336
rect 12671 11308 12716 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 12406 11268 12434 11308
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13357 11339 13415 11345
rect 13357 11305 13369 11339
rect 13403 11336 13415 11339
rect 13814 11336 13820 11348
rect 13403 11308 13820 11336
rect 13403 11305 13415 11308
rect 13357 11299 13415 11305
rect 13814 11296 13820 11308
rect 13872 11336 13878 11348
rect 14274 11336 14280 11348
rect 13872 11308 14280 11336
rect 13872 11296 13878 11308
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 19429 11339 19487 11345
rect 19429 11336 19441 11339
rect 17552 11308 19441 11336
rect 17552 11296 17558 11308
rect 19429 11305 19441 11308
rect 19475 11305 19487 11339
rect 19429 11299 19487 11305
rect 12526 11268 12532 11280
rect 12406 11240 12532 11268
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 17034 11268 17040 11280
rect 14660 11240 17040 11268
rect 3878 11200 3884 11212
rect 1688 11172 3884 11200
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1688 11141 1716 11172
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 5718 11200 5724 11212
rect 4028 11172 5724 11200
rect 4028 11160 4034 11172
rect 5718 11160 5724 11172
rect 5776 11200 5782 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5776 11172 6009 11200
rect 5776 11160 5782 11172
rect 5997 11169 6009 11172
rect 6043 11200 6055 11203
rect 7282 11200 7288 11212
rect 6043 11172 7288 11200
rect 6043 11169 6055 11172
rect 5997 11163 6055 11169
rect 7282 11160 7288 11172
rect 7340 11200 7346 11212
rect 8573 11203 8631 11209
rect 8573 11200 8585 11203
rect 7340 11172 8585 11200
rect 7340 11160 7346 11172
rect 8573 11169 8585 11172
rect 8619 11200 8631 11203
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 8619 11172 9137 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 14660 11200 14688 11240
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 17862 11228 17868 11280
rect 17920 11228 17926 11280
rect 36262 11268 36268 11280
rect 36223 11240 36268 11268
rect 36262 11228 36268 11240
rect 36320 11228 36326 11280
rect 14826 11200 14832 11212
rect 9548 11172 12434 11200
rect 9548 11160 9554 11172
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1636 11104 1685 11132
rect 1636 11092 1642 11104
rect 1673 11101 1685 11104
rect 1719 11101 1731 11135
rect 6546 11132 6552 11144
rect 6507 11104 6552 11132
rect 1673 11095 1731 11101
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11848 11104 11897 11132
rect 11848 11092 11854 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 12406 11132 12434 11172
rect 13280 11172 14688 11200
rect 14787 11172 14832 11200
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 12406 11104 12633 11132
rect 11885 11095 11943 11101
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 13280 11141 13308 11172
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15841 11203 15899 11209
rect 15841 11200 15853 11203
rect 15436 11172 15853 11200
rect 15436 11160 15442 11172
rect 15841 11169 15853 11172
rect 15887 11200 15899 11203
rect 15930 11200 15936 11212
rect 15887 11172 15936 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 16761 11203 16819 11209
rect 16761 11200 16773 11203
rect 16632 11172 16773 11200
rect 16632 11160 16638 11172
rect 16761 11169 16773 11172
rect 16807 11169 16819 11203
rect 16761 11163 16819 11169
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 17880 11200 17908 11228
rect 17451 11172 18644 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 12768 11104 13277 11132
rect 12768 11092 12774 11104
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 1946 11064 1952 11076
rect 1907 11036 1952 11064
rect 1946 11024 1952 11036
rect 2004 11024 2010 11076
rect 3174 11036 4476 11064
rect 4448 10996 4476 11036
rect 4982 11024 4988 11076
rect 5040 11024 5046 11076
rect 5721 11067 5779 11073
rect 5721 11033 5733 11067
rect 5767 11064 5779 11067
rect 6270 11064 6276 11076
rect 5767 11036 6276 11064
rect 5767 11033 5779 11036
rect 5721 11027 5779 11033
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 6822 11024 6828 11076
rect 6880 11024 6886 11076
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 8297 11067 8355 11073
rect 6972 11036 7130 11064
rect 6972 11024 6978 11036
rect 8297 11033 8309 11067
rect 8343 11064 8355 11067
rect 8386 11064 8392 11076
rect 8343 11036 8392 11064
rect 8343 11033 8355 11036
rect 8297 11027 8355 11033
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 9030 11024 9036 11076
rect 9088 11064 9094 11076
rect 9401 11067 9459 11073
rect 9401 11064 9413 11067
rect 9088 11036 9413 11064
rect 9088 11024 9094 11036
rect 9401 11033 9413 11036
rect 9447 11033 9459 11067
rect 9401 11027 9459 11033
rect 9858 11024 9864 11076
rect 9916 11024 9922 11076
rect 11609 11067 11667 11073
rect 11609 11064 11621 11067
rect 10704 11036 11621 11064
rect 5994 10996 6000 11008
rect 4448 10968 6000 10996
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 6840 10996 6868 11024
rect 10704 11008 10732 11036
rect 11609 11033 11621 11036
rect 11655 11033 11667 11067
rect 11609 11027 11667 11033
rect 14369 11067 14427 11073
rect 14369 11033 14381 11067
rect 14415 11033 14427 11067
rect 14369 11027 14427 11033
rect 9214 10996 9220 11008
rect 6840 10968 9220 10996
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 10686 10956 10692 11008
rect 10744 10956 10750 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 14384 10996 14412 11027
rect 14458 11024 14464 11076
rect 14516 11064 14522 11076
rect 14516 11036 14561 11064
rect 14516 11024 14522 11036
rect 14642 11024 14648 11076
rect 14700 11064 14706 11076
rect 16025 11067 16083 11073
rect 16025 11064 16037 11067
rect 14700 11036 16037 11064
rect 14700 11024 14706 11036
rect 16025 11033 16037 11036
rect 16071 11033 16083 11067
rect 16025 11027 16083 11033
rect 16117 11067 16175 11073
rect 16117 11033 16129 11067
rect 16163 11064 16175 11067
rect 16163 11036 16804 11064
rect 16163 11033 16175 11036
rect 16117 11027 16175 11033
rect 15562 10996 15568 11008
rect 12676 10968 15568 10996
rect 12676 10956 12682 10968
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 16776 10996 16804 11036
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 16908 11036 16953 11064
rect 16908 11024 16914 11036
rect 17494 11024 17500 11076
rect 17552 11064 17558 11076
rect 17957 11067 18015 11073
rect 17957 11064 17969 11067
rect 17552 11036 17969 11064
rect 17552 11024 17558 11036
rect 17957 11033 17969 11036
rect 18003 11033 18015 11067
rect 17957 11027 18015 11033
rect 18046 11024 18052 11076
rect 18104 11064 18110 11076
rect 18616 11073 18644 11172
rect 36078 11132 36084 11144
rect 36039 11104 36084 11132
rect 36078 11092 36084 11104
rect 36136 11092 36142 11144
rect 18601 11067 18659 11073
rect 18104 11036 18149 11064
rect 18104 11024 18110 11036
rect 18601 11033 18613 11067
rect 18647 11064 18659 11067
rect 19334 11064 19340 11076
rect 18647 11036 19340 11064
rect 18647 11033 18659 11036
rect 18601 11027 18659 11033
rect 19334 11024 19340 11036
rect 19392 11024 19398 11076
rect 17586 10996 17592 11008
rect 16776 10968 17592 10996
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 1104 10906 36892 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 36892 10906
rect 1104 10832 36892 10854
rect 3878 10792 3884 10804
rect 3839 10764 3884 10792
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 6914 10792 6920 10804
rect 6875 10764 6920 10792
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 7524 10764 10149 10792
rect 7524 10752 7530 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 14550 10792 14556 10804
rect 10137 10755 10195 10761
rect 10244 10764 14556 10792
rect 8478 10684 8484 10736
rect 8536 10684 8542 10736
rect 10244 10724 10272 10764
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 17678 10792 17684 10804
rect 14844 10764 17684 10792
rect 9140 10696 10272 10724
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 2682 10656 2688 10668
rect 2639 10628 2688 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 4985 10619 5043 10625
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 4798 10588 4804 10600
rect 2179 10560 4804 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5000 10520 5028 10619
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 7340 10628 7573 10656
rect 7340 10616 7346 10628
rect 7561 10625 7573 10628
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 7834 10588 7840 10600
rect 7795 10560 7840 10588
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 9140 10588 9168 10696
rect 11698 10684 11704 10736
rect 11756 10724 11762 10736
rect 12253 10727 12311 10733
rect 12253 10724 12265 10727
rect 11756 10696 12265 10724
rect 11756 10684 11762 10696
rect 12253 10693 12265 10696
rect 12299 10693 12311 10727
rect 14090 10724 14096 10736
rect 12253 10687 12311 10693
rect 13096 10696 14096 10724
rect 9214 10616 9220 10668
rect 9272 10656 9278 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 9272 10628 10241 10656
rect 9272 10616 9278 10628
rect 10229 10625 10241 10628
rect 10275 10625 10287 10659
rect 10870 10656 10876 10668
rect 10831 10628 10876 10656
rect 10229 10619 10287 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 13096 10665 13124 10696
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 14734 10724 14740 10736
rect 14695 10696 14740 10724
rect 14734 10684 14740 10696
rect 14792 10684 14798 10736
rect 14844 10733 14872 10764
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 19613 10795 19671 10801
rect 19613 10761 19625 10795
rect 19659 10792 19671 10795
rect 21818 10792 21824 10804
rect 19659 10764 21824 10792
rect 19659 10761 19671 10764
rect 19613 10755 19671 10761
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10693 14887 10727
rect 14829 10687 14887 10693
rect 15838 10684 15844 10736
rect 15896 10724 15902 10736
rect 16025 10727 16083 10733
rect 16025 10724 16037 10727
rect 15896 10696 16037 10724
rect 15896 10684 15902 10696
rect 16025 10693 16037 10696
rect 16071 10693 16083 10727
rect 16025 10687 16083 10693
rect 17037 10727 17095 10733
rect 17037 10693 17049 10727
rect 17083 10724 17095 10727
rect 18506 10724 18512 10736
rect 17083 10696 18512 10724
rect 17083 10693 17095 10696
rect 17037 10687 17095 10693
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13262 10616 13268 10668
rect 13320 10656 13326 10668
rect 13722 10656 13728 10668
rect 13320 10628 13728 10656
rect 13320 10616 13326 10628
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 18877 10659 18935 10665
rect 17644 10628 17689 10656
rect 17644 10616 17650 10628
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 19628 10656 19656 10755
rect 21818 10752 21824 10764
rect 21876 10752 21882 10804
rect 18923 10628 19656 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 9582 10588 9588 10600
rect 8352 10560 9168 10588
rect 9543 10560 9588 10588
rect 8352 10548 8358 10560
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 11606 10548 11612 10600
rect 11664 10588 11670 10600
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11664 10560 11713 10588
rect 11664 10548 11670 10560
rect 11701 10557 11713 10560
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 12345 10591 12403 10597
rect 12345 10557 12357 10591
rect 12391 10588 12403 10591
rect 15654 10588 15660 10600
rect 12391 10560 14412 10588
rect 15615 10560 15660 10588
rect 12391 10557 12403 10560
rect 12345 10551 12403 10557
rect 7558 10520 7564 10532
rect 5000 10492 7564 10520
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 10226 10480 10232 10532
rect 10284 10520 10290 10532
rect 12710 10520 12716 10532
rect 10284 10492 12716 10520
rect 10284 10480 10290 10492
rect 12710 10480 12716 10492
rect 12768 10480 12774 10532
rect 14274 10520 14280 10532
rect 14235 10492 14280 10520
rect 14274 10480 14280 10492
rect 14332 10480 14338 10532
rect 14384 10520 14412 10560
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16942 10588 16948 10600
rect 16163 10560 16948 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 15746 10520 15752 10532
rect 14384 10492 15752 10520
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 4890 10452 4896 10464
rect 4851 10424 4896 10452
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 7282 10452 7288 10464
rect 6043 10424 7288 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 7984 10424 10793 10452
rect 7984 10412 7990 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12032 10424 13001 10452
rect 12032 10412 12038 10424
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 12989 10415 13047 10421
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 13228 10424 13645 10452
rect 13228 10412 13234 10424
rect 13633 10421 13645 10424
rect 13679 10421 13691 10455
rect 14292 10452 14320 10480
rect 14826 10452 14832 10464
rect 14292 10424 14832 10452
rect 13633 10415 13691 10421
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 19061 10455 19119 10461
rect 19061 10421 19073 10455
rect 19107 10452 19119 10455
rect 19426 10452 19432 10464
rect 19107 10424 19432 10452
rect 19107 10421 19119 10424
rect 19061 10415 19119 10421
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 1104 10362 36892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 36892 10362
rect 1104 10288 36892 10310
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4801 10251 4859 10257
rect 4801 10248 4813 10251
rect 4028 10220 4813 10248
rect 4028 10208 4034 10220
rect 4801 10217 4813 10220
rect 4847 10217 4859 10251
rect 8294 10248 8300 10260
rect 4801 10211 4859 10217
rect 5000 10220 8300 10248
rect 3786 10140 3792 10192
rect 3844 10180 3850 10192
rect 4065 10183 4123 10189
rect 4065 10180 4077 10183
rect 3844 10152 4077 10180
rect 3844 10140 3850 10152
rect 4065 10149 4077 10152
rect 4111 10149 4123 10183
rect 4065 10143 4123 10149
rect 1578 10112 1584 10124
rect 1539 10084 1584 10112
rect 1578 10072 1584 10084
rect 1636 10072 1642 10124
rect 1854 10112 1860 10124
rect 1815 10084 1860 10112
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 4614 10112 4620 10124
rect 3375 10084 4620 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 4890 10044 4896 10056
rect 4295 10016 4896 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 5000 10053 5028 10220
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8478 10248 8484 10260
rect 8439 10220 8484 10248
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 15838 10248 15844 10260
rect 11940 10220 12434 10248
rect 15799 10220 15844 10248
rect 11940 10208 11946 10220
rect 7558 10140 7564 10192
rect 7616 10180 7622 10192
rect 10778 10180 10784 10192
rect 7616 10152 10784 10180
rect 7616 10140 7622 10152
rect 10778 10140 10784 10152
rect 10836 10140 10842 10192
rect 12406 10180 12434 10220
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 12713 10183 12771 10189
rect 12713 10180 12725 10183
rect 12406 10152 12725 10180
rect 12713 10149 12725 10152
rect 12759 10149 12771 10183
rect 12713 10143 12771 10149
rect 5718 10112 5724 10124
rect 5679 10084 5724 10112
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 6086 10072 6092 10124
rect 6144 10112 6150 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 6144 10084 9321 10112
rect 6144 10072 6150 10084
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 10594 10112 10600 10124
rect 9309 10075 9367 10081
rect 9416 10084 10600 10112
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 9214 10044 9220 10056
rect 8435 10016 9220 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9416 10053 9444 10084
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10112 11851 10115
rect 11882 10112 11888 10124
rect 11839 10084 11888 10112
rect 11839 10081 11851 10084
rect 11793 10075 11851 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12066 10112 12072 10124
rect 12027 10084 12072 10112
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 13814 10112 13820 10124
rect 13311 10084 13820 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10112 14979 10115
rect 18138 10112 18144 10124
rect 14967 10084 18144 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 10468 10016 11468 10044
rect 10468 10004 10474 10016
rect 5997 9979 6055 9985
rect 3082 9948 5948 9976
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 5258 9908 5264 9920
rect 4856 9880 5264 9908
rect 4856 9868 4862 9880
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 5920 9908 5948 9948
rect 5997 9945 6009 9979
rect 6043 9976 6055 9979
rect 6086 9976 6092 9988
rect 6043 9948 6092 9976
rect 6043 9945 6055 9948
rect 5997 9939 6055 9945
rect 6086 9936 6092 9948
rect 6144 9936 6150 9988
rect 7006 9936 7012 9988
rect 7064 9936 7070 9988
rect 8478 9976 8484 9988
rect 7300 9948 8484 9976
rect 7300 9908 7328 9948
rect 8478 9936 8484 9948
rect 8536 9936 8542 9988
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 10137 9979 10195 9985
rect 10137 9976 10149 9979
rect 9824 9948 10149 9976
rect 9824 9936 9830 9948
rect 10137 9945 10149 9948
rect 10183 9945 10195 9979
rect 11440 9976 11468 10016
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15252 10016 15761 10044
rect 15252 10004 15258 10016
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 11790 9976 11796 9988
rect 10137 9939 10195 9945
rect 10520 9948 11008 9976
rect 11440 9948 11796 9976
rect 7466 9908 7472 9920
rect 5920 9880 7328 9908
rect 7427 9880 7472 9908
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 10520 9908 10548 9948
rect 7892 9880 10548 9908
rect 7892 9868 7898 9880
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 10873 9911 10931 9917
rect 10873 9908 10885 9911
rect 10652 9880 10885 9908
rect 10652 9868 10658 9880
rect 10873 9877 10885 9880
rect 10919 9877 10931 9911
rect 10980 9908 11008 9948
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 11974 9976 11980 9988
rect 11935 9948 11980 9976
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 13170 9976 13176 9988
rect 13131 9948 13176 9976
rect 13170 9936 13176 9948
rect 13228 9936 13234 9988
rect 14274 9976 14280 9988
rect 14235 9948 14280 9976
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 14826 9976 14832 9988
rect 14787 9948 14832 9976
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 14090 9908 14096 9920
rect 10980 9880 14096 9908
rect 10873 9871 10931 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 16482 9908 16488 9920
rect 16443 9880 16488 9908
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 17034 9908 17040 9920
rect 16947 9880 17040 9908
rect 17034 9868 17040 9880
rect 17092 9908 17098 9920
rect 35434 9908 35440 9920
rect 17092 9880 35440 9908
rect 17092 9868 17098 9880
rect 35434 9868 35440 9880
rect 35492 9868 35498 9920
rect 1104 9818 36892 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 36892 9818
rect 1104 9744 36892 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 5534 9704 5540 9716
rect 2740 9676 5540 9704
rect 2740 9664 2746 9676
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 8297 9707 8355 9713
rect 6880 9676 8248 9704
rect 6880 9664 6886 9676
rect 2498 9596 2504 9648
rect 2556 9596 2562 9648
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3142 9636 3148 9648
rect 3099 9608 3148 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3142 9596 3148 9608
rect 3200 9636 3206 9648
rect 3326 9636 3332 9648
rect 3200 9608 3332 9636
rect 3200 9596 3206 9608
rect 3326 9596 3332 9608
rect 3384 9596 3390 9648
rect 5902 9636 5908 9648
rect 5750 9608 5908 9636
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 6972 9608 7314 9636
rect 6972 9596 6978 9608
rect 6546 9568 6552 9580
rect 6507 9540 6552 9568
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 8220 9568 8248 9676
rect 8297 9673 8309 9707
rect 8343 9673 8355 9707
rect 8297 9667 8355 9673
rect 8312 9636 8340 9667
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 9122 9704 9128 9716
rect 8444 9676 9128 9704
rect 8444 9664 8450 9676
rect 9122 9664 9128 9676
rect 9180 9704 9186 9716
rect 9180 9676 9352 9704
rect 9180 9664 9186 9676
rect 8662 9636 8668 9648
rect 8312 9608 8668 9636
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 8754 9568 8760 9580
rect 8220 9540 8760 9568
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 9324 9577 9352 9676
rect 9582 9664 9588 9716
rect 9640 9704 9646 9716
rect 9640 9676 9996 9704
rect 9640 9664 9646 9676
rect 9401 9639 9459 9645
rect 9401 9605 9413 9639
rect 9447 9636 9459 9639
rect 9858 9636 9864 9648
rect 9447 9608 9864 9636
rect 9447 9605 9459 9608
rect 9401 9599 9459 9605
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 9968 9636 9996 9676
rect 12986 9664 12992 9716
rect 13044 9664 13050 9716
rect 16482 9664 16488 9716
rect 16540 9704 16546 9716
rect 17678 9704 17684 9716
rect 16540 9676 17684 9704
rect 16540 9664 16546 9676
rect 17678 9664 17684 9676
rect 17736 9704 17742 9716
rect 36078 9704 36084 9716
rect 17736 9676 36084 9704
rect 17736 9664 17742 9676
rect 36078 9664 36084 9676
rect 36136 9664 36142 9716
rect 9968 9608 11744 9636
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 10229 9571 10287 9577
rect 9355 9540 10180 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 3375 9472 4261 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 4890 9500 4896 9512
rect 4571 9472 4896 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 4264 9364 4292 9463
rect 4890 9460 4896 9472
rect 4948 9500 4954 9512
rect 5166 9500 5172 9512
rect 4948 9472 5172 9500
rect 4948 9460 4954 9472
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 5316 9472 6837 9500
rect 5316 9460 5322 9472
rect 6825 9469 6837 9472
rect 6871 9500 6883 9503
rect 9398 9500 9404 9512
rect 6871 9472 9404 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 10042 9500 10048 9512
rect 9732 9472 10048 9500
rect 9732 9460 9738 9472
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10152 9500 10180 9540
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10318 9568 10324 9580
rect 10275 9540 10324 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10413 9503 10471 9509
rect 10413 9500 10425 9503
rect 10152 9472 10425 9500
rect 10413 9469 10425 9472
rect 10459 9469 10471 9503
rect 11716 9500 11744 9608
rect 12066 9596 12072 9648
rect 12124 9636 12130 9648
rect 12897 9639 12955 9645
rect 12897 9636 12909 9639
rect 12124 9608 12909 9636
rect 12124 9596 12130 9608
rect 12897 9605 12909 9608
rect 12943 9605 12955 9639
rect 13004 9636 13032 9664
rect 14829 9639 14887 9645
rect 13004 9608 13952 9636
rect 12897 9599 12955 9605
rect 11974 9528 11980 9580
rect 12032 9568 12038 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 12032 9540 12173 9568
rect 12032 9528 12038 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9566 13047 9571
rect 13078 9566 13084 9580
rect 13035 9538 13084 9566
rect 13035 9537 13047 9538
rect 12989 9531 13047 9537
rect 13078 9528 13084 9538
rect 13136 9568 13142 9580
rect 13814 9568 13820 9580
rect 13136 9540 13820 9568
rect 13136 9528 13142 9540
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 13924 9577 13952 9608
rect 14829 9605 14841 9639
rect 14875 9636 14887 9639
rect 15010 9636 15016 9648
rect 14875 9608 15016 9636
rect 14875 9605 14887 9608
rect 14829 9599 14887 9605
rect 15010 9596 15016 9608
rect 15068 9596 15074 9648
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9568 13967 9571
rect 14550 9568 14556 9580
rect 13955 9540 14556 9568
rect 13955 9537 13967 9540
rect 13909 9531 13967 9537
rect 14550 9528 14556 9540
rect 14608 9568 14614 9580
rect 14921 9571 14979 9577
rect 14608 9540 14872 9568
rect 14608 9528 14614 9540
rect 12253 9503 12311 9509
rect 11716 9472 12204 9500
rect 10413 9463 10471 9469
rect 6546 9432 6552 9444
rect 5552 9404 6552 9432
rect 5552 9376 5580 9404
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 8846 9432 8852 9444
rect 8128 9404 8852 9432
rect 5534 9364 5540 9376
rect 4264 9336 5540 9364
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5997 9367 6055 9373
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 6086 9364 6092 9376
rect 6043 9336 6092 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 6086 9324 6092 9336
rect 6144 9364 6150 9376
rect 8128 9364 8156 9404
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 10502 9432 10508 9444
rect 9784 9404 10508 9432
rect 6144 9336 8156 9364
rect 6144 9324 6150 9336
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8352 9336 8769 9364
rect 8352 9324 8358 9336
rect 8757 9333 8769 9336
rect 8803 9364 8815 9367
rect 9784 9364 9812 9404
rect 10502 9392 10508 9404
rect 10560 9392 10566 9444
rect 12176 9432 12204 9472
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 14642 9500 14648 9512
rect 12299 9472 14648 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 14844 9500 14872 9540
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 15102 9568 15108 9580
rect 14967 9540 15108 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 18598 9500 18604 9512
rect 14844 9472 18604 9500
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 12986 9432 12992 9444
rect 12176 9404 12992 9432
rect 12986 9392 12992 9404
rect 13044 9392 13050 9444
rect 14274 9432 14280 9444
rect 13096 9404 14280 9432
rect 8803 9336 9812 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 9858 9324 9864 9376
rect 9916 9364 9922 9376
rect 13096 9364 13124 9404
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 9916 9336 13124 9364
rect 9916 9324 9922 9336
rect 13170 9324 13176 9376
rect 13228 9364 13234 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13228 9336 13829 9364
rect 13228 9324 13234 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 15528 9336 15853 9364
rect 15528 9324 15534 9336
rect 15841 9333 15853 9336
rect 15887 9364 15899 9367
rect 27154 9364 27160 9376
rect 15887 9336 27160 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 27154 9324 27160 9336
rect 27212 9324 27218 9376
rect 1104 9274 36892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 36892 9274
rect 1104 9200 36892 9222
rect 3421 9163 3479 9169
rect 3421 9129 3433 9163
rect 3467 9160 3479 9163
rect 3467 9132 5948 9160
rect 3467 9129 3479 9132
rect 3421 9123 3479 9129
rect 5920 9092 5948 9132
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 6549 9163 6607 9169
rect 6549 9160 6561 9163
rect 6052 9132 6561 9160
rect 6052 9120 6058 9132
rect 6549 9129 6561 9132
rect 6595 9129 6607 9163
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 6549 9123 6607 9129
rect 7668 9132 7757 9160
rect 6362 9092 6368 9104
rect 5920 9064 6368 9092
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 7668 9092 7696 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 8478 9160 8484 9172
rect 8439 9132 8484 9160
rect 7745 9123 7803 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 10229 9163 10287 9169
rect 8904 9132 9996 9160
rect 8904 9120 8910 9132
rect 7616 9064 7696 9092
rect 7616 9052 7622 9064
rect 9490 9052 9496 9104
rect 9548 9092 9554 9104
rect 9585 9095 9643 9101
rect 9585 9092 9597 9095
rect 9548 9064 9597 9092
rect 9548 9052 9554 9064
rect 9585 9061 9597 9064
rect 9631 9061 9643 9095
rect 9585 9055 9643 9061
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 5258 9024 5264 9036
rect 4295 8996 5264 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 5997 9027 6055 9033
rect 5997 9024 6009 9027
rect 5776 8996 6009 9024
rect 5776 8984 5782 8996
rect 5997 8993 6009 8996
rect 6043 8993 6055 9027
rect 5997 8987 6055 8993
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 9858 9024 9864 9036
rect 8444 8996 9864 9024
rect 8444 8984 8450 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 9968 9024 9996 9132
rect 10229 9129 10241 9163
rect 10275 9160 10287 9163
rect 11054 9160 11060 9172
rect 10275 9132 11060 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 13265 9163 13323 9169
rect 13265 9129 13277 9163
rect 13311 9160 13323 9163
rect 14826 9160 14832 9172
rect 13311 9132 14832 9160
rect 13311 9129 13323 9132
rect 13265 9123 13323 9129
rect 14826 9120 14832 9132
rect 14884 9120 14890 9172
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 14976 9132 15021 9160
rect 14976 9120 14982 9132
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 10873 9095 10931 9101
rect 10873 9092 10885 9095
rect 10100 9064 10885 9092
rect 10100 9052 10106 9064
rect 10873 9061 10885 9064
rect 10919 9061 10931 9095
rect 10873 9055 10931 9061
rect 12434 9052 12440 9104
rect 12492 9092 12498 9104
rect 14277 9095 14335 9101
rect 14277 9092 14289 9095
rect 12492 9064 14289 9092
rect 12492 9052 12498 9064
rect 14277 9061 14289 9064
rect 14323 9061 14335 9095
rect 36078 9092 36084 9104
rect 36039 9064 36084 9092
rect 14277 9055 14335 9061
rect 36078 9052 36084 9064
rect 36136 9052 36142 9104
rect 12621 9027 12679 9033
rect 9968 8996 12434 9024
rect 4614 8916 4620 8968
rect 4672 8916 4678 8968
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6604 8928 6653 8956
rect 6604 8916 6610 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8956 7343 8959
rect 7466 8956 7472 8968
rect 7331 8928 7472 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7926 8956 7932 8968
rect 7887 8928 7932 8956
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8573 8959 8631 8965
rect 8573 8956 8585 8959
rect 8536 8928 8585 8956
rect 8536 8916 8542 8928
rect 8573 8925 8585 8928
rect 8619 8956 8631 8959
rect 8754 8956 8760 8968
rect 8619 8928 8760 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 9674 8956 9680 8968
rect 9635 8928 9680 8956
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10652 8928 10977 8956
rect 10652 8916 10658 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8925 11943 8959
rect 12406 8956 12434 8996
rect 12621 8993 12633 9027
rect 12667 9024 12679 9027
rect 14734 9024 14740 9036
rect 12667 8996 14740 9024
rect 12667 8993 12679 8996
rect 12621 8987 12679 8993
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12406 8928 12541 8956
rect 11885 8919 11943 8925
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 1946 8888 1952 8900
rect 1907 8860 1952 8888
rect 1946 8848 1952 8860
rect 2004 8848 2010 8900
rect 2038 8848 2044 8900
rect 2096 8888 2102 8900
rect 5721 8891 5779 8897
rect 2096 8860 2438 8888
rect 2096 8848 2102 8860
rect 5721 8857 5733 8891
rect 5767 8857 5779 8891
rect 6086 8888 6092 8900
rect 5721 8851 5779 8857
rect 5920 8860 6092 8888
rect 5736 8820 5764 8851
rect 5920 8820 5948 8860
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 6270 8848 6276 8900
rect 6328 8888 6334 8900
rect 6328 8860 7328 8888
rect 6328 8848 6334 8860
rect 5736 8792 5948 8820
rect 5994 8780 6000 8832
rect 6052 8820 6058 8832
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 6052 8792 7205 8820
rect 6052 8780 6058 8792
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7300 8820 7328 8860
rect 7374 8848 7380 8900
rect 7432 8888 7438 8900
rect 11900 8888 11928 8919
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 12768 8928 13185 8956
rect 12768 8916 12774 8928
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 7432 8860 11928 8888
rect 11977 8891 12035 8897
rect 7432 8848 7438 8860
rect 11977 8857 11989 8891
rect 12023 8888 12035 8891
rect 16850 8888 16856 8900
rect 12023 8860 16856 8888
rect 12023 8857 12035 8860
rect 11977 8851 12035 8857
rect 16850 8848 16856 8860
rect 16908 8848 16914 8900
rect 35621 8891 35679 8897
rect 35621 8857 35633 8891
rect 35667 8888 35679 8891
rect 36262 8888 36268 8900
rect 35667 8860 36268 8888
rect 35667 8857 35679 8860
rect 35621 8851 35679 8857
rect 36262 8848 36268 8860
rect 36320 8848 36326 8900
rect 12526 8820 12532 8832
rect 7300 8792 12532 8820
rect 7193 8783 7251 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 15381 8823 15439 8829
rect 15381 8820 15393 8823
rect 15160 8792 15393 8820
rect 15160 8780 15166 8792
rect 15381 8789 15393 8792
rect 15427 8789 15439 8823
rect 15381 8783 15439 8789
rect 1104 8730 36892 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 36892 8730
rect 1104 8656 36892 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5721 8619 5779 8625
rect 4948 8588 5672 8616
rect 4948 8576 4954 8588
rect 2593 8551 2651 8557
rect 2593 8517 2605 8551
rect 2639 8548 2651 8551
rect 2682 8548 2688 8560
rect 2639 8520 2688 8548
rect 2639 8517 2651 8520
rect 2593 8511 2651 8517
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 3418 8508 3424 8560
rect 3476 8548 3482 8560
rect 3602 8548 3608 8560
rect 3476 8520 3608 8548
rect 3476 8508 3482 8520
rect 3602 8508 3608 8520
rect 3660 8508 3666 8560
rect 4341 8551 4399 8557
rect 4341 8517 4353 8551
rect 4387 8548 4399 8551
rect 5534 8548 5540 8560
rect 4387 8520 5540 8548
rect 4387 8517 4399 8520
rect 4341 8511 4399 8517
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 5644 8548 5672 8588
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5810 8616 5816 8628
rect 5767 8588 5816 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6454 8576 6460 8628
rect 6512 8616 6518 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 6512 8588 7757 8616
rect 6512 8576 6518 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 9306 8616 9312 8628
rect 9267 8588 9312 8616
rect 7745 8579 7803 8585
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11330 8616 11336 8628
rect 11195 8588 11336 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11756 8588 11805 8616
rect 11756 8576 11762 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 11793 8579 11851 8585
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 12805 8619 12863 8625
rect 12805 8616 12817 8619
rect 12492 8588 12817 8616
rect 12492 8576 12498 8588
rect 12805 8585 12817 8588
rect 12851 8616 12863 8619
rect 13446 8616 13452 8628
rect 12851 8588 13452 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 13998 8616 14004 8628
rect 13959 8588 14004 8616
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14550 8616 14556 8628
rect 14511 8588 14556 8616
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 6270 8548 6276 8560
rect 5644 8520 6276 8548
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 7116 8520 8401 8548
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 3878 8480 3884 8492
rect 2179 8452 3884 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4948 8452 4997 8480
rect 4948 8440 4954 8452
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5408 8452 5641 8480
rect 5408 8440 5414 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 7116 8480 7144 8520
rect 8389 8517 8401 8520
rect 8435 8517 8447 8551
rect 9674 8548 9680 8560
rect 8389 8511 8447 8517
rect 9232 8520 9680 8548
rect 6788 8452 7144 8480
rect 7193 8483 7251 8489
rect 6788 8440 6794 8452
rect 7193 8449 7205 8483
rect 7239 8480 7251 8483
rect 7282 8480 7288 8492
rect 7239 8452 7288 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 7208 8412 7236 8443
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7524 8452 7849 8480
rect 7524 8440 7530 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 8478 8480 8484 8492
rect 8439 8452 8484 8480
rect 7837 8443 7895 8449
rect 7742 8412 7748 8424
rect 7208 8384 7748 8412
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 7852 8412 7880 8443
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 9232 8412 9260 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 10134 8548 10140 8560
rect 9876 8520 10140 8548
rect 9398 8480 9404 8492
rect 9359 8452 9404 8480
rect 9398 8440 9404 8452
rect 9456 8480 9462 8492
rect 9876 8480 9904 8520
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 10410 8548 10416 8560
rect 10371 8520 10416 8548
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 10505 8551 10563 8557
rect 10505 8517 10517 8551
rect 10551 8548 10563 8551
rect 11882 8548 11888 8560
rect 10551 8520 11888 8548
rect 10551 8517 10563 8520
rect 10505 8511 10563 8517
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 9456 8452 9904 8480
rect 11701 8483 11759 8489
rect 9456 8440 9462 8452
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 18598 8480 18604 8492
rect 17083 8452 18604 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 7852 8384 9260 8412
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 9861 8415 9919 8421
rect 9861 8412 9873 8415
rect 9364 8384 9873 8412
rect 9364 8372 9370 8384
rect 9861 8381 9873 8384
rect 9907 8412 9919 8415
rect 11606 8412 11612 8424
rect 9907 8384 11612 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 2682 8304 2688 8356
rect 2740 8344 2746 8356
rect 4801 8347 4859 8353
rect 4801 8344 4813 8347
rect 2740 8316 4813 8344
rect 2740 8304 2746 8316
rect 4801 8313 4813 8316
rect 4847 8313 4859 8347
rect 11716 8344 11744 8443
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 4801 8307 4859 8313
rect 4908 8316 11744 8344
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 4908 8276 4936 8316
rect 7098 8276 7104 8288
rect 3476 8248 4936 8276
rect 7059 8248 7104 8276
rect 3476 8236 3482 8248
rect 7098 8236 7104 8248
rect 7156 8236 7162 8288
rect 1104 8186 36892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 36892 8186
rect 1104 8112 36892 8134
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 3418 8072 3424 8084
rect 3292 8044 3424 8072
rect 3292 8032 3298 8044
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 5718 8072 5724 8084
rect 5679 8044 5724 8072
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 7374 8072 7380 8084
rect 6604 8044 7380 8072
rect 6604 8032 6610 8044
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 10962 8072 10968 8084
rect 10919 8044 10968 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 13449 8075 13507 8081
rect 11563 8044 13308 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 5074 7964 5080 8016
rect 5132 8004 5138 8016
rect 7469 8007 7527 8013
rect 7469 8004 7481 8007
rect 5132 7976 7481 8004
rect 5132 7964 5138 7976
rect 7469 7973 7481 7976
rect 7515 7973 7527 8007
rect 13078 8004 13084 8016
rect 7469 7967 7527 7973
rect 12406 7976 13084 8004
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 4249 7939 4307 7945
rect 1995 7908 3832 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 3050 7828 3056 7880
rect 3108 7828 3114 7880
rect 3804 7812 3832 7908
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 4295 7908 7236 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 5684 7840 7021 7868
rect 5684 7828 5690 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7208 7868 7236 7908
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7340 7908 11468 7936
rect 7340 7896 7346 7908
rect 8294 7868 8300 7880
rect 7208 7840 8300 7868
rect 7009 7831 7067 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8573 7871 8631 7877
rect 8573 7868 8585 7871
rect 8536 7840 8585 7868
rect 8536 7828 8542 7840
rect 8573 7837 8585 7840
rect 8619 7868 8631 7871
rect 8938 7868 8944 7880
rect 8619 7840 8944 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 11440 7877 11468 7908
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9272 7840 9413 7868
rect 9272 7828 9278 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 10781 7871 10839 7877
rect 10781 7868 10793 7871
rect 9401 7831 9459 7837
rect 9508 7840 10793 7868
rect 3786 7760 3792 7812
rect 3844 7800 3850 7812
rect 9508 7800 9536 7840
rect 10781 7837 10793 7840
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 3844 7772 9536 7800
rect 9677 7803 9735 7809
rect 3844 7760 3850 7772
rect 9677 7769 9689 7803
rect 9723 7769 9735 7803
rect 9677 7763 9735 7769
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 5500 7704 8493 7732
rect 5500 7692 5506 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 8481 7695 8539 7701
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 9692 7732 9720 7763
rect 8996 7704 9720 7732
rect 8996 7692 9002 7704
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 12161 7735 12219 7741
rect 12161 7732 12173 7735
rect 12032 7704 12173 7732
rect 12032 7692 12038 7704
rect 12161 7701 12173 7704
rect 12207 7732 12219 7735
rect 12406 7732 12434 7976
rect 13078 7964 13084 7976
rect 13136 7964 13142 8016
rect 13280 8004 13308 8044
rect 13449 8041 13461 8075
rect 13495 8072 13507 8075
rect 13722 8072 13728 8084
rect 13495 8044 13728 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 36173 8075 36231 8081
rect 36173 8041 36185 8075
rect 36219 8072 36231 8075
rect 36630 8072 36636 8084
rect 36219 8044 36636 8072
rect 36219 8041 36231 8044
rect 36173 8035 36231 8041
rect 36630 8032 36636 8044
rect 36688 8032 36694 8084
rect 14182 8004 14188 8016
rect 13280 7976 14188 8004
rect 14182 7964 14188 7976
rect 14240 7964 14246 8016
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7936 12863 7939
rect 14090 7936 14096 7948
rect 12851 7908 14096 7936
rect 12851 7905 12863 7908
rect 12805 7899 12863 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 35621 7803 35679 7809
rect 35621 7769 35633 7803
rect 35667 7800 35679 7803
rect 36262 7800 36268 7812
rect 35667 7772 36268 7800
rect 35667 7769 35679 7772
rect 35621 7763 35679 7769
rect 36262 7760 36268 7772
rect 36320 7760 36326 7812
rect 12207 7704 12434 7732
rect 12207 7701 12219 7704
rect 12161 7695 12219 7701
rect 1104 7642 36892 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 36892 7642
rect 1104 7568 36892 7590
rect 3786 7528 3792 7540
rect 3747 7500 3792 7528
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 5534 7528 5540 7540
rect 3988 7500 5540 7528
rect 2590 7420 2596 7472
rect 2648 7420 2654 7472
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 3142 7460 3148 7472
rect 2832 7432 3148 7460
rect 2832 7420 2838 7432
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7392 3387 7395
rect 3418 7392 3424 7404
rect 3375 7364 3424 7392
rect 3375 7361 3387 7364
rect 3329 7355 3387 7361
rect 3418 7352 3424 7364
rect 3476 7392 3482 7404
rect 3988 7392 4016 7500
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 6638 7528 6644 7540
rect 6599 7500 6644 7528
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7837 7531 7895 7537
rect 7837 7497 7849 7531
rect 7883 7528 7895 7531
rect 8110 7528 8116 7540
rect 7883 7500 8116 7528
rect 7883 7497 7895 7500
rect 7837 7491 7895 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8389 7531 8447 7537
rect 8389 7497 8401 7531
rect 8435 7528 8447 7531
rect 10410 7528 10416 7540
rect 8435 7500 10416 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12437 7531 12495 7537
rect 12437 7528 12449 7531
rect 12308 7500 12449 7528
rect 12308 7488 12314 7500
rect 12437 7497 12449 7500
rect 12483 7497 12495 7531
rect 12437 7491 12495 7497
rect 5258 7460 5264 7472
rect 4830 7432 5264 7460
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 9582 7460 9588 7472
rect 5736 7432 9588 7460
rect 3476 7364 4016 7392
rect 3476 7352 3482 7364
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5592 7364 5637 7392
rect 5592 7352 5598 7364
rect 5736 7336 5764 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 6546 7392 6552 7404
rect 6507 7364 6552 7392
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 8297 7395 8355 7401
rect 8297 7392 8309 7395
rect 6656 7364 8309 7392
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7324 3111 7327
rect 5166 7324 5172 7336
rect 3099 7296 5172 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7324 5319 7327
rect 5718 7324 5724 7336
rect 5307 7296 5724 7324
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 1946 7256 1952 7268
rect 1627 7228 1952 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 1946 7216 1952 7228
rect 2004 7216 2010 7268
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 6656 7188 6684 7364
rect 8297 7361 8309 7364
rect 8343 7361 8355 7395
rect 9214 7392 9220 7404
rect 9127 7364 9220 7392
rect 8297 7355 8355 7361
rect 9214 7352 9220 7364
rect 9272 7392 9278 7404
rect 9766 7392 9772 7404
rect 9272 7364 9772 7392
rect 9272 7352 9278 7364
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12986 7392 12992 7404
rect 12023 7364 12992 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 9398 7324 9404 7336
rect 9359 7296 9404 7324
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 7285 7259 7343 7265
rect 7285 7225 7297 7259
rect 7331 7256 7343 7259
rect 9674 7256 9680 7268
rect 7331 7228 9680 7256
rect 7331 7225 7343 7228
rect 7285 7219 7343 7225
rect 9674 7216 9680 7228
rect 9732 7256 9738 7268
rect 10594 7256 10600 7268
rect 9732 7228 10600 7256
rect 9732 7216 9738 7228
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 3752 7160 6684 7188
rect 3752 7148 3758 7160
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10318 7188 10324 7200
rect 9824 7160 10324 7188
rect 9824 7148 9830 7160
rect 10318 7148 10324 7160
rect 10376 7188 10382 7200
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 10376 7160 11805 7188
rect 10376 7148 10382 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 11793 7151 11851 7157
rect 1104 7098 36892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 36892 7098
rect 1104 7024 36892 7046
rect 1936 6987 1994 6993
rect 1936 6953 1948 6987
rect 1982 6984 1994 6987
rect 8662 6984 8668 6996
rect 1982 6956 8668 6984
rect 1982 6953 1994 6956
rect 1936 6947 1994 6953
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 1670 6848 1676 6860
rect 1583 6820 1676 6848
rect 1670 6808 1676 6820
rect 1728 6848 1734 6860
rect 3418 6848 3424 6860
rect 1728 6820 3424 6848
rect 1728 6808 1734 6820
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 5258 6848 5264 6860
rect 5219 6820 5264 6848
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5902 6848 5908 6860
rect 5863 6820 5908 6848
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 7466 6848 7472 6860
rect 7427 6820 7472 6848
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 8570 6848 8576 6860
rect 8531 6820 8576 6848
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 10226 6808 10232 6860
rect 10284 6848 10290 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 10284 6820 10333 6848
rect 10284 6808 10290 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 10594 6808 10600 6860
rect 10652 6848 10658 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 10652 6820 11069 6848
rect 10652 6808 10658 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4709 6783 4767 6789
rect 4709 6780 4721 6783
rect 3844 6752 4721 6780
rect 3844 6740 3850 6752
rect 4709 6749 4721 6752
rect 4755 6749 4767 6783
rect 5350 6780 5356 6792
rect 5311 6752 5356 6780
rect 4709 6743 4767 6749
rect 5350 6740 5356 6752
rect 5408 6780 5414 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5408 6752 6009 6780
rect 5408 6740 5414 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 2958 6672 2964 6724
rect 3016 6672 3022 6724
rect 4617 6715 4675 6721
rect 4617 6712 4629 6715
rect 3344 6684 4629 6712
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 3344 6644 3372 6684
rect 4617 6681 4629 6684
rect 4663 6681 4675 6715
rect 6012 6712 6040 6743
rect 6178 6740 6184 6792
rect 6236 6780 6242 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 6236 6752 9137 6780
rect 6236 6740 6242 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 22373 6783 22431 6789
rect 22373 6780 22385 6783
rect 19392 6752 22385 6780
rect 19392 6740 19398 6752
rect 22373 6749 22385 6752
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 9398 6712 9404 6724
rect 6012 6684 9404 6712
rect 4617 6675 4675 6681
rect 9398 6672 9404 6684
rect 9456 6672 9462 6724
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 12621 6715 12679 6721
rect 12621 6712 12633 6715
rect 11940 6684 12633 6712
rect 11940 6672 11946 6684
rect 12621 6681 12633 6684
rect 12667 6681 12679 6715
rect 13170 6712 13176 6724
rect 13131 6684 13176 6712
rect 12621 6675 12679 6681
rect 13170 6672 13176 6684
rect 13228 6672 13234 6724
rect 13262 6672 13268 6724
rect 13320 6712 13326 6724
rect 13320 6684 13365 6712
rect 13320 6672 13326 6684
rect 2648 6616 3372 6644
rect 3421 6647 3479 6653
rect 2648 6604 2654 6616
rect 3421 6613 3433 6647
rect 3467 6644 3479 6647
rect 3602 6644 3608 6656
rect 3467 6616 3608 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 7009 6647 7067 6653
rect 7009 6613 7021 6647
rect 7055 6644 7067 6647
rect 7650 6644 7656 6656
rect 7055 6616 7656 6644
rect 7055 6613 7067 6616
rect 7009 6607 7067 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 8202 6604 8208 6656
rect 8260 6644 8266 6656
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 8260 6616 9689 6644
rect 8260 6604 8266 6616
rect 9677 6613 9689 6616
rect 9723 6644 9735 6647
rect 17218 6644 17224 6656
rect 9723 6616 17224 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 22465 6647 22523 6653
rect 22465 6613 22477 6647
rect 22511 6644 22523 6647
rect 24670 6644 24676 6656
rect 22511 6616 24676 6644
rect 22511 6613 22523 6616
rect 22465 6607 22523 6613
rect 24670 6604 24676 6616
rect 24728 6604 24734 6656
rect 1104 6554 36892 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 36892 6554
rect 1104 6480 36892 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 3694 6440 3700 6452
rect 1719 6412 3700 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 4249 6443 4307 6449
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 4614 6440 4620 6452
rect 4295 6412 4620 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5684 6412 5917 6440
rect 5684 6400 5690 6412
rect 5905 6409 5917 6412
rect 5951 6440 5963 6443
rect 6546 6440 6552 6452
rect 5951 6412 6552 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 7469 6443 7527 6449
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 7834 6440 7840 6452
rect 7515 6412 7840 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 7834 6400 7840 6412
rect 7892 6400 7898 6452
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7984 6412 8033 6440
rect 7984 6400 7990 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 9030 6440 9036 6452
rect 8991 6412 9036 6440
rect 8021 6403 8079 6409
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9585 6443 9643 6449
rect 9585 6409 9597 6443
rect 9631 6440 9643 6443
rect 9674 6440 9680 6452
rect 9631 6412 9680 6440
rect 9631 6409 9643 6412
rect 9585 6403 9643 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 12989 6443 13047 6449
rect 12989 6409 13001 6443
rect 13035 6440 13047 6443
rect 13262 6440 13268 6452
rect 13035 6412 13268 6440
rect 13035 6409 13047 6412
rect 12989 6403 13047 6409
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 36170 6440 36176 6452
rect 17276 6412 36176 6440
rect 17276 6400 17282 6412
rect 36170 6400 36176 6412
rect 36228 6400 36234 6452
rect 3145 6375 3203 6381
rect 3145 6341 3157 6375
rect 3191 6372 3203 6375
rect 3234 6372 3240 6384
rect 3191 6344 3240 6372
rect 3191 6341 3203 6344
rect 3145 6335 3203 6341
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 4893 6375 4951 6381
rect 4893 6341 4905 6375
rect 4939 6372 4951 6375
rect 7006 6372 7012 6384
rect 4939 6344 7012 6372
rect 4939 6341 4951 6344
rect 4893 6335 4951 6341
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 7742 6332 7748 6384
rect 7800 6372 7806 6384
rect 10045 6375 10103 6381
rect 10045 6372 10057 6375
rect 7800 6344 10057 6372
rect 7800 6332 7806 6344
rect 10045 6341 10057 6344
rect 10091 6341 10103 6375
rect 10045 6335 10103 6341
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 3476 6276 3521 6304
rect 3476 6264 3482 6276
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4157 6307 4215 6313
rect 4157 6304 4169 6307
rect 4120 6276 4169 6304
rect 4120 6264 4126 6276
rect 4157 6273 4169 6276
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 5350 6304 5356 6316
rect 4847 6276 5356 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 4816 6236 4844 6267
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 22094 6304 22100 6316
rect 22055 6276 22100 6304
rect 22094 6264 22100 6276
rect 22152 6304 22158 6316
rect 22741 6307 22799 6313
rect 22741 6304 22753 6307
rect 22152 6276 22753 6304
rect 22152 6264 22158 6276
rect 22741 6273 22753 6276
rect 22787 6273 22799 6307
rect 22741 6267 22799 6273
rect 2648 6208 4844 6236
rect 2648 6196 2654 6208
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 8478 6168 8484 6180
rect 4120 6140 8484 6168
rect 4120 6128 4126 6140
rect 8478 6128 8484 6140
rect 8536 6128 8542 6180
rect 22281 6171 22339 6177
rect 22281 6137 22293 6171
rect 22327 6168 22339 6171
rect 24578 6168 24584 6180
rect 22327 6140 24584 6168
rect 22327 6137 22339 6140
rect 22281 6131 22339 6137
rect 24578 6128 24584 6140
rect 24636 6128 24642 6180
rect 1104 6010 36892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 36892 6010
rect 1104 5936 36892 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 1762 5896 1768 5908
rect 1719 5868 1768 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 1762 5856 1768 5868
rect 1820 5856 1826 5908
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2924 5868 2973 5896
rect 2924 5856 2930 5868
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 2961 5859 3019 5865
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3200 5868 4077 5896
rect 3200 5856 3206 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5169 5899 5227 5905
rect 5169 5896 5181 5899
rect 4856 5868 5181 5896
rect 4856 5856 4862 5868
rect 5169 5865 5181 5868
rect 5215 5865 5227 5899
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 5169 5859 5227 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 6604 5868 7849 5896
rect 6604 5856 6610 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 6641 5831 6699 5837
rect 6641 5828 6653 5831
rect 3844 5800 6653 5828
rect 3844 5788 3850 5800
rect 6641 5797 6653 5800
rect 6687 5828 6699 5831
rect 7285 5831 7343 5837
rect 7285 5828 7297 5831
rect 6687 5800 7297 5828
rect 6687 5797 6699 5800
rect 6641 5791 6699 5797
rect 7285 5797 7297 5800
rect 7331 5828 7343 5831
rect 7742 5828 7748 5840
rect 7331 5800 7748 5828
rect 7331 5797 7343 5800
rect 7285 5791 7343 5797
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 9766 5760 9772 5772
rect 1780 5732 2774 5760
rect 1780 5701 1808 5732
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 2406 5692 2412 5704
rect 2367 5664 2412 5692
rect 1765 5655 1823 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 2746 5692 2774 5732
rect 3068 5732 9772 5760
rect 3068 5701 3096 5732
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2746 5664 3065 5692
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 3234 5652 3240 5704
rect 3292 5692 3298 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3292 5664 3985 5692
rect 3292 5652 3298 5664
rect 3973 5661 3985 5664
rect 4019 5692 4031 5695
rect 4062 5692 4068 5704
rect 4019 5664 4068 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 36081 5695 36139 5701
rect 36081 5692 36093 5695
rect 35866 5664 36093 5692
rect 2314 5624 2320 5636
rect 2275 5596 2320 5624
rect 2314 5584 2320 5596
rect 2372 5584 2378 5636
rect 3602 5584 3608 5636
rect 3660 5624 3666 5636
rect 4617 5627 4675 5633
rect 4617 5624 4629 5627
rect 3660 5596 4629 5624
rect 3660 5584 3666 5596
rect 4617 5593 4629 5596
rect 4663 5624 4675 5627
rect 12250 5624 12256 5636
rect 4663 5596 12256 5624
rect 4663 5593 4675 5596
rect 4617 5587 4675 5593
rect 12250 5584 12256 5596
rect 12308 5584 12314 5636
rect 35526 5624 35532 5636
rect 35487 5596 35532 5624
rect 35526 5584 35532 5596
rect 35584 5624 35590 5636
rect 35866 5624 35894 5664
rect 36081 5661 36093 5664
rect 36127 5661 36139 5695
rect 36081 5655 36139 5661
rect 35584 5596 35894 5624
rect 35584 5584 35590 5596
rect 36262 5556 36268 5568
rect 36223 5528 36268 5556
rect 36262 5516 36268 5528
rect 36320 5516 36326 5568
rect 1104 5466 36892 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 36892 5466
rect 1104 5392 36892 5414
rect 2685 5355 2743 5361
rect 2685 5321 2697 5355
rect 2731 5352 2743 5355
rect 3050 5352 3056 5364
rect 2731 5324 3056 5352
rect 2731 5321 2743 5324
rect 2685 5315 2743 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 4706 5352 4712 5364
rect 4663 5324 4712 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5626 5352 5632 5364
rect 5215 5324 5632 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 17678 5352 17684 5364
rect 5776 5324 5821 5352
rect 17639 5324 17684 5352
rect 5776 5312 5782 5324
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 2406 5244 2412 5296
rect 2464 5284 2470 5296
rect 2464 5256 4108 5284
rect 2464 5244 2470 5256
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 1872 5148 1900 5179
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2590 5216 2596 5228
rect 2004 5188 2596 5216
rect 2004 5176 2010 5188
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 4080 5225 4108 5256
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17696 5216 17724 5312
rect 16991 5188 17724 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 5994 5148 6000 5160
rect 1872 5120 6000 5148
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 3329 5083 3387 5089
rect 3329 5049 3341 5083
rect 3375 5080 3387 5083
rect 6914 5080 6920 5092
rect 3375 5052 6920 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 1670 5012 1676 5024
rect 1631 4984 1676 5012
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 3878 5012 3884 5024
rect 3839 4984 3884 5012
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 17129 5015 17187 5021
rect 17129 4981 17141 5015
rect 17175 5012 17187 5015
rect 17494 5012 17500 5024
rect 17175 4984 17500 5012
rect 17175 4981 17187 4984
rect 17129 4975 17187 4981
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 1104 4922 36892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 36892 4922
rect 1104 4848 36892 4870
rect 2038 4808 2044 4820
rect 1999 4780 2044 4808
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 2685 4811 2743 4817
rect 2685 4777 2697 4811
rect 2731 4808 2743 4811
rect 2958 4808 2964 4820
rect 2731 4780 2964 4808
rect 2731 4777 2743 4780
rect 2685 4771 2743 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3326 4808 3332 4820
rect 3287 4780 3332 4808
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3568 4780 3985 4808
rect 3568 4768 3574 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 3973 4771 4031 4777
rect 4709 4811 4767 4817
rect 4709 4777 4721 4811
rect 4755 4808 4767 4811
rect 4890 4808 4896 4820
rect 4755 4780 4896 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5626 4808 5632 4820
rect 5307 4780 5632 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 1946 4604 1952 4616
rect 1907 4576 1952 4604
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 3234 4604 3240 4616
rect 2823 4576 3240 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 9306 4604 9312 4616
rect 9267 4576 9312 4604
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 36078 4604 36084 4616
rect 36039 4576 36084 4604
rect 36078 4564 36084 4576
rect 36136 4564 36142 4616
rect 9214 4468 9220 4480
rect 9175 4440 9220 4468
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 36262 4468 36268 4480
rect 36223 4440 36268 4468
rect 36262 4428 36268 4440
rect 36320 4428 36326 4480
rect 1104 4378 36892 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 36892 4378
rect 1104 4304 36892 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2593 4267 2651 4273
rect 2593 4264 2605 4267
rect 2464 4236 2605 4264
rect 2464 4224 2470 4236
rect 2593 4233 2605 4236
rect 2639 4233 2651 4267
rect 2593 4227 2651 4233
rect 3145 4267 3203 4273
rect 3145 4233 3157 4267
rect 3191 4264 3203 4267
rect 3786 4264 3792 4276
rect 3191 4236 3792 4264
rect 3191 4233 3203 4236
rect 3145 4227 3203 4233
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2774 4128 2780 4140
rect 2455 4100 2780 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 3970 4128 3976 4140
rect 3927 4100 3976 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 25682 4088 25688 4140
rect 25740 4128 25746 4140
rect 25869 4131 25927 4137
rect 25869 4128 25881 4131
rect 25740 4100 25881 4128
rect 25740 4088 25746 4100
rect 25869 4097 25881 4100
rect 25915 4128 25927 4131
rect 26513 4131 26571 4137
rect 26513 4128 26525 4131
rect 25915 4100 26525 4128
rect 25915 4097 25927 4100
rect 25869 4091 25927 4097
rect 26513 4097 26525 4100
rect 26559 4097 26571 4131
rect 26513 4091 26571 4097
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 4982 4060 4988 4072
rect 1903 4032 4988 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 26053 3995 26111 4001
rect 26053 3961 26065 3995
rect 26099 3992 26111 3995
rect 26099 3964 26234 3992
rect 26099 3961 26111 3964
rect 26053 3955 26111 3961
rect 26206 3924 26234 3964
rect 36078 3924 36084 3936
rect 26206 3896 36084 3924
rect 36078 3884 36084 3896
rect 36136 3884 36142 3936
rect 1104 3834 36892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 36892 3834
rect 1104 3760 36892 3782
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 2774 3720 2780 3732
rect 2455 3692 2780 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 3878 3516 3884 3528
rect 1903 3488 3884 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 15988 3488 19441 3516
rect 15988 3476 15994 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 35621 3519 35679 3525
rect 35621 3485 35633 3519
rect 35667 3516 35679 3519
rect 35802 3516 35808 3528
rect 35667 3488 35808 3516
rect 35667 3485 35679 3488
rect 35621 3479 35679 3485
rect 35802 3476 35808 3488
rect 35860 3516 35866 3528
rect 36265 3519 36323 3525
rect 36265 3516 36277 3519
rect 35860 3488 36277 3516
rect 35860 3476 35866 3488
rect 36265 3485 36277 3488
rect 36311 3485 36323 3519
rect 36265 3479 36323 3485
rect 20346 3408 20352 3460
rect 20404 3448 20410 3460
rect 36081 3451 36139 3457
rect 36081 3448 36093 3451
rect 20404 3420 36093 3448
rect 20404 3408 20410 3420
rect 36081 3417 36093 3420
rect 36127 3417 36139 3451
rect 36081 3411 36139 3417
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 19521 3383 19579 3389
rect 19521 3349 19533 3383
rect 19567 3380 19579 3383
rect 20714 3380 20720 3392
rect 19567 3352 20720 3380
rect 19567 3349 19579 3352
rect 19521 3343 19579 3349
rect 20714 3340 20720 3352
rect 20772 3340 20778 3392
rect 1104 3290 36892 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 36892 3290
rect 1104 3216 36892 3238
rect 35434 3176 35440 3188
rect 35395 3148 35440 3176
rect 35434 3136 35440 3148
rect 35492 3136 35498 3188
rect 36170 3176 36176 3188
rect 36131 3148 36176 3176
rect 36170 3136 36176 3148
rect 36228 3136 36234 3188
rect 36722 3108 36728 3120
rect 35866 3080 36728 3108
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 7282 3040 7288 3052
rect 1903 3012 2452 3040
rect 7243 3012 7288 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2424 2913 2452 3012
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 34885 3043 34943 3049
rect 34885 3009 34897 3043
rect 34931 3040 34943 3043
rect 35529 3043 35587 3049
rect 35529 3040 35541 3043
rect 34931 3012 35541 3040
rect 34931 3009 34943 3012
rect 34885 3003 34943 3009
rect 35529 3009 35541 3012
rect 35575 3040 35587 3043
rect 35866 3040 35894 3080
rect 36722 3068 36728 3080
rect 36780 3068 36786 3120
rect 35575 3012 35894 3040
rect 36265 3043 36323 3049
rect 35575 3009 35587 3012
rect 35529 3003 35587 3009
rect 36265 3009 36277 3043
rect 36311 3040 36323 3043
rect 36354 3040 36360 3052
rect 36311 3012 36360 3040
rect 36311 3009 36323 3012
rect 36265 3003 36323 3009
rect 36354 3000 36360 3012
rect 36412 3000 36418 3052
rect 18874 2972 18880 2984
rect 2746 2944 18880 2972
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2904 2467 2907
rect 2746 2904 2774 2944
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 2455 2876 2774 2904
rect 2455 2873 2467 2876
rect 2409 2867 2467 2873
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 7469 2839 7527 2845
rect 7469 2805 7481 2839
rect 7515 2836 7527 2839
rect 7834 2836 7840 2848
rect 7515 2808 7840 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 18785 2839 18843 2845
rect 18785 2805 18797 2839
rect 18831 2836 18843 2839
rect 20622 2836 20628 2848
rect 18831 2808 20628 2836
rect 18831 2805 18843 2808
rect 18785 2799 18843 2805
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 27062 2796 27068 2848
rect 27120 2836 27126 2848
rect 27157 2839 27215 2845
rect 27157 2836 27169 2839
rect 27120 2808 27169 2836
rect 27120 2796 27126 2808
rect 27157 2805 27169 2808
rect 27203 2805 27215 2839
rect 30374 2836 30380 2848
rect 30335 2808 30380 2836
rect 27157 2799 27215 2805
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 1104 2746 36892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 36892 2746
rect 1104 2672 36892 2694
rect 4203 2635 4261 2641
rect 4203 2601 4215 2635
rect 4249 2632 4261 2635
rect 7282 2632 7288 2644
rect 4249 2604 7288 2632
rect 4249 2601 4261 2604
rect 4203 2595 4261 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 12986 2632 12992 2644
rect 12947 2604 12992 2632
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 18598 2632 18604 2644
rect 14507 2604 18604 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 29822 2632 29828 2644
rect 29783 2604 29828 2632
rect 29822 2592 29828 2604
rect 29880 2592 29886 2644
rect 30558 2632 30564 2644
rect 30519 2604 30564 2632
rect 30558 2592 30564 2604
rect 30616 2592 30622 2644
rect 32398 2632 32404 2644
rect 32359 2604 32404 2632
rect 32398 2592 32404 2604
rect 32456 2592 32462 2644
rect 33778 2592 33784 2644
rect 33836 2632 33842 2644
rect 34977 2635 35035 2641
rect 34977 2632 34989 2635
rect 33836 2604 34989 2632
rect 33836 2592 33842 2604
rect 34977 2601 34989 2604
rect 35023 2601 35035 2635
rect 34977 2595 35035 2601
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 72 2536 2421 2564
rect 72 2524 78 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 11974 2564 11980 2576
rect 11935 2536 11980 2564
rect 2409 2527 2467 2533
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 16301 2567 16359 2573
rect 16301 2533 16313 2567
rect 16347 2564 16359 2567
rect 19058 2564 19064 2576
rect 16347 2536 19064 2564
rect 16347 2533 16359 2536
rect 16301 2527 16359 2533
rect 19058 2524 19064 2536
rect 19116 2524 19122 2576
rect 23658 2564 23664 2576
rect 20088 2536 23664 2564
rect 7558 2496 7564 2508
rect 1872 2468 7564 2496
rect 1872 2437 1900 2468
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 20088 2496 20116 2536
rect 23658 2524 23664 2536
rect 23716 2524 23722 2576
rect 27154 2564 27160 2576
rect 27115 2536 27160 2564
rect 27154 2524 27160 2536
rect 27212 2524 27218 2576
rect 33873 2567 33931 2573
rect 33873 2533 33885 2567
rect 33919 2564 33931 2567
rect 34514 2564 34520 2576
rect 33919 2536 34520 2564
rect 33919 2533 33931 2536
rect 33873 2527 33931 2533
rect 34514 2524 34520 2536
rect 34572 2524 34578 2576
rect 7668 2468 20116 2496
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2682 2428 2688 2440
rect 2639 2400 2688 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3344 2400 3985 2428
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3344 2301 3372 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 6871 2400 7389 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 7377 2397 7389 2400
rect 7423 2428 7435 2431
rect 7668 2428 7696 2468
rect 20622 2456 20628 2508
rect 20680 2496 20686 2508
rect 20680 2468 22692 2496
rect 20680 2456 20686 2468
rect 7834 2428 7840 2440
rect 7423 2400 7696 2428
rect 7795 2400 7840 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 5552 2360 5580 2391
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10091 2400 12848 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 9214 2360 9220 2372
rect 5552 2332 9220 2360
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 9309 2363 9367 2369
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 9674 2360 9680 2372
rect 9355 2332 9680 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 9674 2320 9680 2332
rect 9732 2360 9738 2372
rect 9861 2363 9919 2369
rect 9861 2360 9873 2363
rect 9732 2332 9873 2360
rect 9732 2320 9738 2332
rect 9861 2329 9873 2332
rect 9907 2329 9919 2363
rect 9861 2323 9919 2329
rect 11793 2363 11851 2369
rect 11793 2329 11805 2363
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 4580 2264 5365 2292
rect 4580 2252 4586 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 11054 2292 11060 2304
rect 11015 2264 11060 2292
rect 8021 2255 8079 2261
rect 11054 2252 11060 2264
rect 11112 2292 11118 2304
rect 11808 2292 11836 2323
rect 11112 2264 11836 2292
rect 12820 2292 12848 2400
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12952 2400 13185 2428
rect 12952 2388 12958 2400
rect 13173 2397 13185 2400
rect 13219 2428 13231 2431
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13219 2400 13645 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14240 2400 14289 2428
rect 14240 2388 14246 2400
rect 14277 2397 14289 2400
rect 14323 2428 14335 2431
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14323 2400 14933 2428
rect 14323 2397 14335 2400
rect 14277 2391 14335 2397
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 14921 2391 14979 2397
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 20714 2428 20720 2440
rect 20675 2400 20720 2428
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 22664 2437 22692 2468
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 24578 2428 24584 2440
rect 24539 2400 24584 2428
rect 22649 2391 22707 2397
rect 24578 2388 24584 2400
rect 24636 2388 24642 2440
rect 24670 2388 24676 2440
rect 24728 2428 24734 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 24728 2400 25881 2428
rect 24728 2388 24734 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 30432 2400 30665 2428
rect 30432 2388 30438 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 34992 2428 35020 2595
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 34992 2400 35541 2428
rect 30653 2391 30711 2397
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 16114 2360 16120 2372
rect 16075 2332 16120 2360
rect 16114 2320 16120 2332
rect 16172 2360 16178 2372
rect 16853 2363 16911 2369
rect 16853 2360 16865 2363
rect 16172 2332 16865 2360
rect 16172 2320 16178 2332
rect 16853 2329 16865 2332
rect 16899 2329 16911 2363
rect 25682 2360 25688 2372
rect 16853 2323 16911 2329
rect 17328 2332 25688 2360
rect 15102 2292 15108 2304
rect 12820 2264 15108 2292
rect 11112 2252 11118 2264
rect 15102 2252 15108 2264
rect 15160 2292 15166 2304
rect 17328 2292 17356 2332
rect 25682 2320 25688 2332
rect 25740 2320 25746 2372
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27341 2363 27399 2369
rect 27341 2360 27353 2363
rect 27120 2332 27353 2360
rect 27120 2320 27126 2332
rect 27341 2329 27353 2332
rect 27387 2329 27399 2363
rect 29917 2363 29975 2369
rect 29917 2360 29929 2363
rect 27341 2323 27399 2329
rect 29104 2332 29929 2360
rect 15160 2264 17356 2292
rect 15160 2252 15166 2264
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 22833 2255 22891 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24765 2295 24823 2301
rect 24765 2292 24777 2295
rect 23900 2264 24777 2292
rect 23900 2252 23906 2264
rect 24765 2261 24777 2264
rect 24811 2261 24823 2295
rect 24765 2255 24823 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 29104 2301 29132 2332
rect 29917 2329 29929 2332
rect 29963 2329 29975 2363
rect 29917 2323 29975 2329
rect 31757 2363 31815 2369
rect 31757 2329 31769 2363
rect 31803 2360 31815 2363
rect 32214 2360 32220 2372
rect 31803 2332 32220 2360
rect 31803 2329 31815 2332
rect 31757 2323 31815 2329
rect 32214 2320 32220 2332
rect 32272 2360 32278 2372
rect 32493 2363 32551 2369
rect 32493 2360 32505 2363
rect 32272 2332 32505 2360
rect 32272 2320 32278 2332
rect 32493 2329 32505 2332
rect 32539 2329 32551 2363
rect 32493 2323 32551 2329
rect 33137 2363 33195 2369
rect 33137 2329 33149 2363
rect 33183 2360 33195 2363
rect 33502 2360 33508 2372
rect 33183 2332 33508 2360
rect 33183 2329 33195 2332
rect 33137 2323 33195 2329
rect 33502 2320 33508 2332
rect 33560 2360 33566 2372
rect 33689 2363 33747 2369
rect 33689 2360 33701 2363
rect 33560 2332 33701 2360
rect 33560 2320 33566 2332
rect 33689 2329 33701 2332
rect 33735 2329 33747 2363
rect 33689 2323 33747 2329
rect 29089 2295 29147 2301
rect 29089 2292 29101 2295
rect 29052 2264 29101 2292
rect 29052 2252 29058 2264
rect 29089 2261 29101 2264
rect 29135 2261 29147 2295
rect 29089 2255 29147 2261
rect 35434 2252 35440 2304
rect 35492 2292 35498 2304
rect 35713 2295 35771 2301
rect 35713 2292 35725 2295
rect 35492 2264 35725 2292
rect 35492 2252 35498 2264
rect 35713 2261 35725 2264
rect 35759 2261 35771 2295
rect 36354 2292 36360 2304
rect 36315 2264 36360 2292
rect 35713 2255 35771 2261
rect 36354 2252 36360 2264
rect 36412 2252 36418 2304
rect 1104 2202 36892 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 36892 2202
rect 1104 2128 36892 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 14832 37408 14884 37460
rect 26424 37408 26476 37460
rect 2320 37247 2372 37256
rect 2320 37213 2329 37247
rect 2329 37213 2363 37247
rect 2363 37213 2372 37247
rect 2320 37204 2372 37213
rect 3240 37204 3292 37256
rect 4252 37247 4304 37256
rect 4252 37213 4261 37247
rect 4261 37213 4295 37247
rect 4295 37213 4304 37247
rect 4252 37204 4304 37213
rect 5172 37204 5224 37256
rect 7104 37272 7156 37324
rect 16120 37272 16172 37324
rect 26424 37272 26476 37324
rect 32864 37408 32916 37460
rect 34152 37408 34204 37460
rect 32956 37315 33008 37324
rect 32956 37281 32965 37315
rect 32965 37281 32999 37315
rect 32999 37281 33008 37315
rect 32956 37272 33008 37281
rect 9404 37247 9456 37256
rect 9404 37213 9413 37247
rect 9413 37213 9447 37247
rect 9447 37213 9456 37247
rect 9404 37204 9456 37213
rect 10692 37247 10744 37256
rect 10692 37213 10701 37247
rect 10701 37213 10735 37247
rect 10735 37213 10744 37247
rect 10692 37204 10744 37213
rect 10784 37204 10836 37256
rect 14004 37204 14056 37256
rect 14832 37204 14884 37256
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 18052 37204 18104 37256
rect 18880 37204 18932 37256
rect 22008 37247 22060 37256
rect 22008 37213 22017 37247
rect 22017 37213 22051 37247
rect 22051 37213 22060 37247
rect 22008 37204 22060 37213
rect 23296 37247 23348 37256
rect 23296 37213 23305 37247
rect 23305 37213 23339 37247
rect 23339 37213 23348 37247
rect 23296 37204 23348 37213
rect 24584 37247 24636 37256
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 27436 37247 27488 37256
rect 27436 37213 27445 37247
rect 27445 37213 27479 37247
rect 27479 37213 27488 37247
rect 27436 37204 27488 37213
rect 28448 37247 28500 37256
rect 28448 37213 28457 37247
rect 28457 37213 28491 37247
rect 28491 37213 28500 37247
rect 28448 37204 28500 37213
rect 29092 37204 29144 37256
rect 31024 37247 31076 37256
rect 31024 37213 31033 37247
rect 31033 37213 31067 37247
rect 31067 37213 31076 37247
rect 31024 37204 31076 37213
rect 34796 37272 34848 37324
rect 35624 37204 35676 37256
rect 2964 37136 3016 37188
rect 1952 37068 2004 37120
rect 2872 37111 2924 37120
rect 2872 37077 2881 37111
rect 2881 37077 2915 37111
rect 2915 37077 2924 37111
rect 2872 37068 2924 37077
rect 3884 37068 3936 37120
rect 8392 37068 8444 37120
rect 10324 37068 10376 37120
rect 11612 37068 11664 37120
rect 13544 37111 13596 37120
rect 13544 37077 13553 37111
rect 13553 37077 13587 37111
rect 13587 37077 13596 37111
rect 13544 37068 13596 37077
rect 15016 37111 15068 37120
rect 15016 37077 15025 37111
rect 15025 37077 15059 37111
rect 15059 37077 15068 37111
rect 15016 37068 15068 37077
rect 16764 37068 16816 37120
rect 18144 37111 18196 37120
rect 18144 37077 18153 37111
rect 18153 37077 18187 37111
rect 18187 37077 18196 37111
rect 18144 37068 18196 37077
rect 19984 37068 20036 37120
rect 21272 37068 21324 37120
rect 23204 37068 23256 37120
rect 24492 37068 24544 37120
rect 27712 37068 27764 37120
rect 29644 37068 29696 37120
rect 30932 37068 30984 37120
rect 36084 37068 36136 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4252 36864 4304 36916
rect 1676 36839 1728 36848
rect 1676 36805 1685 36839
rect 1685 36805 1719 36839
rect 1719 36805 1728 36839
rect 1676 36796 1728 36805
rect 10692 36864 10744 36916
rect 28448 36864 28500 36916
rect 29092 36907 29144 36916
rect 29092 36873 29101 36907
rect 29101 36873 29135 36907
rect 29135 36873 29144 36907
rect 29092 36864 29144 36873
rect 35532 36907 35584 36916
rect 12256 36796 12308 36848
rect 27436 36796 27488 36848
rect 10876 36728 10928 36780
rect 18144 36728 18196 36780
rect 27160 36771 27212 36780
rect 27160 36737 27169 36771
rect 27169 36737 27203 36771
rect 27203 36737 27212 36771
rect 27160 36728 27212 36737
rect 1860 36635 1912 36644
rect 1860 36601 1869 36635
rect 1869 36601 1903 36635
rect 1903 36601 1912 36635
rect 1860 36592 1912 36601
rect 35532 36873 35541 36907
rect 35541 36873 35575 36907
rect 35575 36873 35584 36907
rect 35532 36864 35584 36873
rect 37372 36796 37424 36848
rect 3240 36567 3292 36576
rect 3240 36533 3249 36567
rect 3249 36533 3283 36567
rect 3283 36533 3292 36567
rect 3240 36524 3292 36533
rect 14004 36524 14056 36576
rect 28356 36567 28408 36576
rect 28356 36533 28365 36567
rect 28365 36533 28399 36567
rect 28399 36533 28408 36567
rect 28356 36524 28408 36533
rect 36176 36567 36228 36576
rect 36176 36533 36185 36567
rect 36185 36533 36219 36567
rect 36219 36533 36228 36567
rect 36176 36524 36228 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 17684 36320 17736 36372
rect 28356 36320 28408 36372
rect 35624 36363 35676 36372
rect 35624 36329 35633 36363
rect 35633 36329 35667 36363
rect 35667 36329 35676 36363
rect 35624 36320 35676 36329
rect 2504 36252 2556 36304
rect 664 36116 716 36168
rect 26424 36116 26476 36168
rect 36268 36023 36320 36032
rect 36268 35989 36277 36023
rect 36277 35989 36311 36023
rect 36311 35989 36320 36023
rect 36268 35980 36320 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1584 35615 1636 35624
rect 1584 35581 1593 35615
rect 1593 35581 1627 35615
rect 1627 35581 1636 35615
rect 1584 35572 1636 35581
rect 2688 35572 2740 35624
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1584 35275 1636 35284
rect 1584 35241 1593 35275
rect 1593 35241 1627 35275
rect 1627 35241 1636 35275
rect 1584 35232 1636 35241
rect 27160 35028 27212 35080
rect 36360 35071 36412 35080
rect 36360 35037 36369 35071
rect 36369 35037 36403 35071
rect 36403 35037 36412 35071
rect 36360 35028 36412 35037
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 36360 34731 36412 34740
rect 36360 34697 36369 34731
rect 36369 34697 36403 34731
rect 36403 34697 36412 34731
rect 36360 34688 36412 34697
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 18880 33099 18932 33108
rect 18880 33065 18889 33099
rect 18889 33065 18923 33099
rect 18923 33065 18932 33099
rect 18880 33056 18932 33065
rect 18236 32852 18288 32904
rect 13820 32784 13872 32836
rect 31024 32784 31076 32836
rect 36268 32827 36320 32836
rect 36268 32793 36277 32827
rect 36277 32793 36311 32827
rect 36311 32793 36320 32827
rect 36268 32784 36320 32793
rect 36544 32716 36596 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1584 32351 1636 32360
rect 1584 32317 1593 32351
rect 1593 32317 1627 32351
rect 1627 32317 1636 32351
rect 1584 32308 1636 32317
rect 2780 32308 2832 32360
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1584 32011 1636 32020
rect 1584 31977 1593 32011
rect 1593 31977 1627 32011
rect 1627 31977 1636 32011
rect 1584 31968 1636 31977
rect 10784 31968 10836 32020
rect 35808 31900 35860 31952
rect 5724 31764 5776 31816
rect 10692 31807 10744 31816
rect 10692 31773 10701 31807
rect 10701 31773 10735 31807
rect 10735 31773 10744 31807
rect 10692 31764 10744 31773
rect 10876 31764 10928 31816
rect 27804 31764 27856 31816
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 9404 31424 9456 31476
rect 12900 31288 12952 31340
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 24584 30880 24636 30932
rect 13176 30676 13228 30728
rect 21180 30676 21232 30728
rect 1676 30583 1728 30592
rect 1676 30549 1685 30583
rect 1685 30549 1719 30583
rect 1719 30549 1728 30583
rect 1676 30540 1728 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 13176 30379 13228 30388
rect 13176 30345 13185 30379
rect 13185 30345 13219 30379
rect 13219 30345 13228 30379
rect 13176 30336 13228 30345
rect 2320 30268 2372 30320
rect 4620 30200 4672 30252
rect 12532 30200 12584 30252
rect 12624 30200 12676 30252
rect 12256 30107 12308 30116
rect 12256 30073 12265 30107
rect 12265 30073 12299 30107
rect 12299 30073 12308 30107
rect 12256 30064 12308 30073
rect 27436 30200 27488 30252
rect 32956 30064 33008 30116
rect 22560 30039 22612 30048
rect 22560 30005 22569 30039
rect 22569 30005 22603 30039
rect 22603 30005 22612 30039
rect 22560 29996 22612 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 27160 29588 27212 29640
rect 36268 29563 36320 29572
rect 36268 29529 36277 29563
rect 36277 29529 36311 29563
rect 36311 29529 36320 29563
rect 36268 29520 36320 29529
rect 12532 29495 12584 29504
rect 12532 29461 12541 29495
rect 12541 29461 12575 29495
rect 12575 29461 12584 29495
rect 12532 29452 12584 29461
rect 17224 29452 17276 29504
rect 35992 29452 36044 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 16120 29291 16172 29300
rect 16120 29257 16129 29291
rect 16129 29257 16163 29291
rect 16163 29257 16172 29291
rect 16120 29248 16172 29257
rect 1584 29155 1636 29164
rect 1584 29121 1593 29155
rect 1593 29121 1627 29155
rect 1627 29121 1636 29155
rect 1584 29112 1636 29121
rect 1768 29019 1820 29028
rect 1768 28985 1777 29019
rect 1777 28985 1811 29019
rect 1811 28985 1820 29019
rect 1768 28976 1820 28985
rect 15660 28976 15712 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 16856 28704 16908 28756
rect 13912 28500 13964 28552
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 36268 28067 36320 28076
rect 36268 28033 36277 28067
rect 36277 28033 36311 28067
rect 36311 28033 36320 28067
rect 36268 28024 36320 28033
rect 15568 27888 15620 27940
rect 35900 27888 35952 27940
rect 1860 27820 1912 27872
rect 12072 27820 12124 27872
rect 15476 27820 15528 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 12624 27591 12676 27600
rect 12624 27557 12633 27591
rect 12633 27557 12667 27591
rect 12667 27557 12676 27591
rect 12624 27548 12676 27557
rect 1860 27455 1912 27464
rect 1860 27421 1869 27455
rect 1869 27421 1903 27455
rect 1903 27421 1912 27455
rect 1860 27412 1912 27421
rect 2504 27455 2556 27464
rect 2504 27421 2513 27455
rect 2513 27421 2547 27455
rect 2547 27421 2556 27455
rect 2504 27412 2556 27421
rect 15476 27412 15528 27464
rect 2688 27344 2740 27396
rect 16396 27344 16448 27396
rect 1676 27319 1728 27328
rect 1676 27285 1685 27319
rect 1685 27285 1719 27319
rect 1719 27285 1728 27319
rect 1676 27276 1728 27285
rect 2320 27319 2372 27328
rect 2320 27285 2329 27319
rect 2329 27285 2363 27319
rect 2363 27285 2372 27319
rect 2320 27276 2372 27285
rect 11152 27276 11204 27328
rect 11796 27276 11848 27328
rect 14464 27276 14516 27328
rect 14832 27319 14884 27328
rect 14832 27285 14841 27319
rect 14841 27285 14875 27319
rect 14875 27285 14884 27319
rect 14832 27276 14884 27285
rect 14924 27276 14976 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 5908 27072 5960 27124
rect 8576 27004 8628 27056
rect 11796 27047 11848 27056
rect 11796 27013 11805 27047
rect 11805 27013 11839 27047
rect 11839 27013 11848 27047
rect 11796 27004 11848 27013
rect 11888 27047 11940 27056
rect 11888 27013 11897 27047
rect 11897 27013 11931 27047
rect 11931 27013 11940 27047
rect 11888 27004 11940 27013
rect 13820 27004 13872 27056
rect 14188 27004 14240 27056
rect 14924 27047 14976 27056
rect 14924 27013 14933 27047
rect 14933 27013 14967 27047
rect 14967 27013 14976 27047
rect 14924 27004 14976 27013
rect 15660 27047 15712 27056
rect 15660 27013 15669 27047
rect 15669 27013 15703 27047
rect 15703 27013 15712 27047
rect 15660 27004 15712 27013
rect 16672 27004 16724 27056
rect 2964 26936 3016 26988
rect 11152 26979 11204 26988
rect 11152 26945 11161 26979
rect 11161 26945 11195 26979
rect 11195 26945 11204 26979
rect 11152 26936 11204 26945
rect 16396 26936 16448 26988
rect 7932 26911 7984 26920
rect 7932 26877 7941 26911
rect 7941 26877 7975 26911
rect 7975 26877 7984 26911
rect 7932 26868 7984 26877
rect 12072 26868 12124 26920
rect 1492 26800 1544 26852
rect 4988 26800 5040 26852
rect 9220 26800 9272 26852
rect 10600 26800 10652 26852
rect 15844 26868 15896 26920
rect 17592 26868 17644 26920
rect 1952 26732 2004 26784
rect 10508 26775 10560 26784
rect 10508 26741 10517 26775
rect 10517 26741 10551 26775
rect 10551 26741 10560 26775
rect 10508 26732 10560 26741
rect 10968 26732 11020 26784
rect 16580 26732 16632 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 6736 26528 6788 26580
rect 1860 26460 1912 26512
rect 8208 26460 8260 26512
rect 10600 26460 10652 26512
rect 5264 26392 5316 26444
rect 7932 26435 7984 26444
rect 7932 26401 7941 26435
rect 7941 26401 7975 26435
rect 7975 26401 7984 26435
rect 7932 26392 7984 26401
rect 9220 26435 9272 26444
rect 9220 26401 9229 26435
rect 9229 26401 9263 26435
rect 9263 26401 9272 26435
rect 9220 26392 9272 26401
rect 10692 26392 10744 26444
rect 11888 26528 11940 26580
rect 12440 26460 12492 26512
rect 1676 26324 1728 26376
rect 3608 26324 3660 26376
rect 12256 26324 12308 26376
rect 12624 26324 12676 26376
rect 2688 26256 2740 26308
rect 9772 26299 9824 26308
rect 9772 26265 9781 26299
rect 9781 26265 9815 26299
rect 9815 26265 9824 26299
rect 9772 26256 9824 26265
rect 10968 26299 11020 26308
rect 10968 26265 10977 26299
rect 10977 26265 11011 26299
rect 11011 26265 11020 26299
rect 10968 26256 11020 26265
rect 12900 26435 12952 26444
rect 12900 26401 12909 26435
rect 12909 26401 12943 26435
rect 12943 26401 12952 26435
rect 12900 26392 12952 26401
rect 15844 26392 15896 26444
rect 17224 26528 17276 26580
rect 17500 26460 17552 26512
rect 35808 26460 35860 26512
rect 17316 26435 17368 26444
rect 17316 26401 17325 26435
rect 17325 26401 17359 26435
rect 17359 26401 17368 26435
rect 17316 26392 17368 26401
rect 22560 26392 22612 26444
rect 14556 26324 14608 26376
rect 15292 26324 15344 26376
rect 36084 26367 36136 26376
rect 36084 26333 36093 26367
rect 36093 26333 36127 26367
rect 36127 26333 36136 26367
rect 36084 26324 36136 26333
rect 15384 26299 15436 26308
rect 15384 26265 15393 26299
rect 15393 26265 15427 26299
rect 15427 26265 15436 26299
rect 15384 26256 15436 26265
rect 14372 26188 14424 26240
rect 17592 26256 17644 26308
rect 18512 26256 18564 26308
rect 16856 26188 16908 26240
rect 16948 26188 17000 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 3240 25984 3292 26036
rect 8300 25984 8352 26036
rect 8576 26027 8628 26036
rect 8576 25993 8585 26027
rect 8585 25993 8619 26027
rect 8619 25993 8628 26027
rect 8576 25984 8628 25993
rect 9772 25984 9824 26036
rect 2136 25959 2188 25968
rect 2136 25925 2145 25959
rect 2145 25925 2179 25959
rect 2179 25925 2188 25959
rect 2136 25916 2188 25925
rect 2504 25916 2556 25968
rect 5264 25959 5316 25968
rect 2596 25848 2648 25900
rect 5264 25925 5273 25959
rect 5273 25925 5307 25959
rect 5307 25925 5316 25959
rect 5264 25916 5316 25925
rect 9680 25916 9732 25968
rect 10692 25916 10744 25968
rect 15016 25984 15068 26036
rect 13268 25959 13320 25968
rect 13268 25925 13277 25959
rect 13277 25925 13311 25959
rect 13311 25925 13320 25959
rect 13268 25916 13320 25925
rect 14372 25959 14424 25968
rect 14372 25925 14381 25959
rect 14381 25925 14415 25959
rect 14415 25925 14424 25959
rect 14372 25916 14424 25925
rect 17500 25984 17552 26036
rect 17040 25916 17092 25968
rect 8760 25848 8812 25900
rect 9220 25891 9272 25900
rect 9220 25857 9229 25891
rect 9229 25857 9263 25891
rect 9263 25857 9272 25891
rect 9220 25848 9272 25857
rect 12072 25891 12124 25900
rect 2044 25780 2096 25832
rect 2504 25780 2556 25832
rect 2688 25780 2740 25832
rect 4988 25780 5040 25832
rect 10140 25780 10192 25832
rect 10508 25780 10560 25832
rect 12072 25857 12081 25891
rect 12081 25857 12115 25891
rect 12115 25857 12124 25891
rect 12072 25848 12124 25857
rect 15568 25891 15620 25900
rect 15568 25857 15577 25891
rect 15577 25857 15611 25891
rect 15611 25857 15620 25891
rect 15568 25848 15620 25857
rect 18236 25891 18288 25900
rect 12716 25823 12768 25832
rect 12716 25789 12725 25823
rect 12725 25789 12759 25823
rect 12759 25789 12768 25823
rect 12716 25780 12768 25789
rect 13360 25823 13412 25832
rect 13360 25789 13369 25823
rect 13369 25789 13403 25823
rect 13403 25789 13412 25823
rect 13360 25780 13412 25789
rect 5724 25755 5776 25764
rect 3516 25687 3568 25696
rect 3516 25653 3525 25687
rect 3525 25653 3559 25687
rect 3559 25653 3568 25687
rect 3516 25644 3568 25653
rect 5724 25721 5733 25755
rect 5733 25721 5767 25755
rect 5767 25721 5776 25755
rect 5724 25712 5776 25721
rect 11336 25712 11388 25764
rect 15292 25780 15344 25832
rect 18236 25857 18245 25891
rect 18245 25857 18279 25891
rect 18279 25857 18288 25891
rect 18236 25848 18288 25857
rect 35900 25848 35952 25900
rect 16580 25780 16632 25832
rect 17224 25780 17276 25832
rect 17500 25823 17552 25832
rect 17500 25789 17509 25823
rect 17509 25789 17543 25823
rect 17543 25789 17552 25823
rect 17500 25780 17552 25789
rect 16212 25712 16264 25764
rect 6828 25644 6880 25696
rect 7932 25687 7984 25696
rect 7932 25653 7941 25687
rect 7941 25653 7975 25687
rect 7975 25653 7984 25687
rect 7932 25644 7984 25653
rect 10508 25644 10560 25696
rect 11244 25644 11296 25696
rect 12164 25687 12216 25696
rect 12164 25653 12173 25687
rect 12173 25653 12207 25687
rect 12207 25653 12216 25687
rect 12164 25644 12216 25653
rect 13820 25644 13872 25696
rect 17776 25644 17828 25696
rect 18144 25687 18196 25696
rect 18144 25653 18153 25687
rect 18153 25653 18187 25687
rect 18187 25653 18196 25687
rect 18144 25644 18196 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3516 25440 3568 25492
rect 12532 25440 12584 25492
rect 14740 25440 14792 25492
rect 16212 25440 16264 25492
rect 17040 25483 17092 25492
rect 17040 25449 17049 25483
rect 17049 25449 17083 25483
rect 17083 25449 17092 25483
rect 17040 25440 17092 25449
rect 2044 25304 2096 25356
rect 4620 25372 4672 25424
rect 8208 25372 8260 25424
rect 8300 25372 8352 25424
rect 2412 25211 2464 25220
rect 2412 25177 2421 25211
rect 2421 25177 2455 25211
rect 2455 25177 2464 25211
rect 2412 25168 2464 25177
rect 10968 25347 11020 25356
rect 10968 25313 10977 25347
rect 10977 25313 11011 25347
rect 11011 25313 11020 25347
rect 10968 25304 11020 25313
rect 11336 25347 11388 25356
rect 11336 25313 11345 25347
rect 11345 25313 11379 25347
rect 11379 25313 11388 25347
rect 11336 25304 11388 25313
rect 12164 25304 12216 25356
rect 13360 25372 13412 25424
rect 20076 25440 20128 25492
rect 17868 25372 17920 25424
rect 18144 25304 18196 25356
rect 22560 25304 22612 25356
rect 3332 25279 3384 25288
rect 3332 25245 3341 25279
rect 3341 25245 3375 25279
rect 3375 25245 3384 25279
rect 3332 25236 3384 25245
rect 5540 25236 5592 25288
rect 9680 25236 9732 25288
rect 9956 25279 10008 25288
rect 9956 25245 9965 25279
rect 9965 25245 9999 25279
rect 9999 25245 10008 25279
rect 9956 25236 10008 25245
rect 3792 25168 3844 25220
rect 5816 25211 5868 25220
rect 5816 25177 5825 25211
rect 5825 25177 5859 25211
rect 5859 25177 5868 25211
rect 5816 25168 5868 25177
rect 3148 25143 3200 25152
rect 3148 25109 3157 25143
rect 3157 25109 3191 25143
rect 3191 25109 3200 25143
rect 3148 25100 3200 25109
rect 4436 25100 4488 25152
rect 4988 25100 5040 25152
rect 5172 25143 5224 25152
rect 5172 25109 5181 25143
rect 5181 25109 5215 25143
rect 5215 25109 5224 25143
rect 5172 25100 5224 25109
rect 5448 25100 5500 25152
rect 7012 25211 7064 25220
rect 7012 25177 7021 25211
rect 7021 25177 7055 25211
rect 7055 25177 7064 25211
rect 7012 25168 7064 25177
rect 8208 25168 8260 25220
rect 9496 25168 9548 25220
rect 11244 25211 11296 25220
rect 11244 25177 11253 25211
rect 11253 25177 11287 25211
rect 11287 25177 11296 25211
rect 11244 25168 11296 25177
rect 8852 25100 8904 25152
rect 9864 25143 9916 25152
rect 9864 25109 9873 25143
rect 9873 25109 9907 25143
rect 9907 25109 9916 25143
rect 9864 25100 9916 25109
rect 10600 25100 10652 25152
rect 11612 25168 11664 25220
rect 12256 25168 12308 25220
rect 13636 25279 13688 25288
rect 13636 25245 13645 25279
rect 13645 25245 13679 25279
rect 13679 25245 13688 25279
rect 13636 25236 13688 25245
rect 14832 25236 14884 25288
rect 16488 25236 16540 25288
rect 14096 25168 14148 25220
rect 14464 25211 14516 25220
rect 14464 25177 14473 25211
rect 14473 25177 14507 25211
rect 14507 25177 14516 25211
rect 14464 25168 14516 25177
rect 15476 25168 15528 25220
rect 15292 25143 15344 25152
rect 15292 25109 15301 25143
rect 15301 25109 15335 25143
rect 15335 25109 15344 25143
rect 15292 25100 15344 25109
rect 16028 25143 16080 25152
rect 16028 25109 16037 25143
rect 16037 25109 16071 25143
rect 16071 25109 16080 25143
rect 16028 25100 16080 25109
rect 17776 25211 17828 25220
rect 17776 25177 17785 25211
rect 17785 25177 17819 25211
rect 17819 25177 17828 25211
rect 20812 25211 20864 25220
rect 17776 25168 17828 25177
rect 20812 25177 20821 25211
rect 20821 25177 20855 25211
rect 20855 25177 20864 25211
rect 20812 25168 20864 25177
rect 18052 25100 18104 25152
rect 18788 25143 18840 25152
rect 18788 25109 18797 25143
rect 18797 25109 18831 25143
rect 18831 25109 18840 25143
rect 18788 25100 18840 25109
rect 19248 25100 19300 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 2228 24828 2280 24880
rect 1952 24692 2004 24744
rect 3792 24828 3844 24880
rect 3884 24871 3936 24880
rect 3884 24837 3893 24871
rect 3893 24837 3927 24871
rect 3927 24837 3936 24871
rect 3884 24828 3936 24837
rect 5540 24828 5592 24880
rect 6644 24828 6696 24880
rect 7288 24828 7340 24880
rect 7932 24828 7984 24880
rect 10508 24871 10560 24880
rect 2780 24803 2832 24812
rect 2780 24769 2789 24803
rect 2789 24769 2823 24803
rect 2823 24769 2832 24803
rect 2780 24760 2832 24769
rect 5632 24760 5684 24812
rect 5908 24803 5960 24812
rect 5908 24769 5917 24803
rect 5917 24769 5951 24803
rect 5951 24769 5960 24803
rect 5908 24760 5960 24769
rect 7380 24803 7432 24812
rect 4528 24624 4580 24676
rect 4436 24556 4488 24608
rect 4988 24692 5040 24744
rect 7380 24769 7389 24803
rect 7389 24769 7423 24803
rect 7423 24769 7432 24803
rect 7380 24760 7432 24769
rect 8116 24760 8168 24812
rect 8668 24803 8720 24812
rect 8668 24769 8677 24803
rect 8677 24769 8711 24803
rect 8711 24769 8720 24803
rect 10508 24837 10517 24871
rect 10517 24837 10551 24871
rect 10551 24837 10560 24871
rect 10508 24828 10560 24837
rect 10968 24896 11020 24948
rect 15384 24896 15436 24948
rect 16028 24896 16080 24948
rect 33784 24896 33836 24948
rect 11612 24828 11664 24880
rect 11888 24871 11940 24880
rect 11888 24837 11897 24871
rect 11897 24837 11931 24871
rect 11931 24837 11940 24871
rect 11888 24828 11940 24837
rect 13544 24828 13596 24880
rect 14832 24871 14884 24880
rect 14832 24837 14841 24871
rect 14841 24837 14875 24871
rect 14875 24837 14884 24871
rect 14832 24828 14884 24837
rect 17040 24871 17092 24880
rect 17040 24837 17049 24871
rect 17049 24837 17083 24871
rect 17083 24837 17092 24871
rect 17040 24828 17092 24837
rect 17132 24828 17184 24880
rect 17776 24828 17828 24880
rect 8668 24760 8720 24769
rect 9956 24760 10008 24812
rect 14188 24803 14240 24812
rect 14188 24769 14197 24803
rect 14197 24769 14231 24803
rect 14231 24769 14240 24803
rect 18512 24803 18564 24812
rect 14188 24760 14240 24769
rect 18512 24769 18521 24803
rect 18521 24769 18555 24803
rect 18555 24769 18564 24803
rect 18512 24760 18564 24769
rect 18604 24803 18656 24812
rect 18604 24769 18613 24803
rect 18613 24769 18647 24803
rect 18647 24769 18656 24803
rect 18604 24760 18656 24769
rect 18788 24760 18840 24812
rect 21088 24760 21140 24812
rect 6736 24692 6788 24744
rect 6184 24624 6236 24676
rect 6368 24624 6420 24676
rect 8668 24624 8720 24676
rect 4804 24556 4856 24608
rect 4896 24556 4948 24608
rect 8024 24556 8076 24608
rect 8944 24556 8996 24608
rect 10048 24667 10100 24676
rect 10048 24633 10057 24667
rect 10057 24633 10091 24667
rect 10091 24633 10100 24667
rect 10600 24735 10652 24744
rect 10600 24701 10609 24735
rect 10609 24701 10643 24735
rect 10643 24701 10652 24735
rect 10600 24692 10652 24701
rect 11336 24692 11388 24744
rect 13268 24692 13320 24744
rect 13360 24692 13412 24744
rect 14740 24735 14792 24744
rect 14740 24701 14749 24735
rect 14749 24701 14783 24735
rect 14783 24701 14792 24735
rect 14740 24692 14792 24701
rect 12348 24667 12400 24676
rect 10048 24624 10100 24633
rect 12348 24633 12357 24667
rect 12357 24633 12391 24667
rect 12391 24633 12400 24667
rect 12348 24624 12400 24633
rect 14464 24624 14516 24676
rect 17132 24692 17184 24744
rect 17316 24692 17368 24744
rect 35900 24692 35952 24744
rect 36360 24735 36412 24744
rect 36360 24701 36369 24735
rect 36369 24701 36403 24735
rect 36403 24701 36412 24735
rect 36360 24692 36412 24701
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 17316 24556 17368 24608
rect 19248 24556 19300 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2136 24352 2188 24404
rect 3332 24352 3384 24404
rect 5816 24352 5868 24404
rect 7012 24395 7064 24404
rect 7012 24361 7021 24395
rect 7021 24361 7055 24395
rect 7055 24361 7064 24395
rect 7012 24352 7064 24361
rect 7104 24352 7156 24404
rect 1400 24284 1452 24336
rect 1768 24216 1820 24268
rect 1952 24148 2004 24200
rect 4896 24216 4948 24268
rect 5264 24216 5316 24268
rect 5080 24148 5132 24200
rect 6736 24148 6788 24200
rect 7104 24191 7156 24200
rect 7104 24157 7113 24191
rect 7113 24157 7147 24191
rect 7147 24157 7156 24191
rect 7104 24148 7156 24157
rect 7840 24191 7892 24200
rect 7840 24157 7849 24191
rect 7849 24157 7883 24191
rect 7883 24157 7892 24191
rect 9220 24284 9272 24336
rect 13544 24352 13596 24404
rect 15568 24352 15620 24404
rect 20812 24352 20864 24404
rect 36360 24395 36412 24404
rect 36360 24361 36369 24395
rect 36369 24361 36403 24395
rect 36403 24361 36412 24395
rect 36360 24352 36412 24361
rect 12716 24284 12768 24336
rect 12992 24284 13044 24336
rect 13728 24284 13780 24336
rect 14740 24284 14792 24336
rect 9496 24259 9548 24268
rect 9496 24225 9505 24259
rect 9505 24225 9539 24259
rect 9539 24225 9548 24259
rect 9496 24216 9548 24225
rect 11060 24216 11112 24268
rect 12164 24259 12216 24268
rect 12164 24225 12173 24259
rect 12173 24225 12207 24259
rect 12207 24225 12216 24259
rect 12164 24216 12216 24225
rect 12440 24259 12492 24268
rect 12440 24225 12449 24259
rect 12449 24225 12483 24259
rect 12483 24225 12492 24259
rect 12440 24216 12492 24225
rect 12808 24216 12860 24268
rect 13176 24216 13228 24268
rect 14188 24216 14240 24268
rect 16488 24216 16540 24268
rect 17500 24216 17552 24268
rect 18144 24216 18196 24268
rect 7840 24148 7892 24157
rect 17224 24148 17276 24200
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 4620 24055 4672 24064
rect 4620 24021 4629 24055
rect 4629 24021 4663 24055
rect 4663 24021 4672 24055
rect 4620 24012 4672 24021
rect 5356 24012 5408 24064
rect 8484 24012 8536 24064
rect 10784 24123 10836 24132
rect 10784 24089 10793 24123
rect 10793 24089 10827 24123
rect 10827 24089 10836 24123
rect 10784 24080 10836 24089
rect 10048 24012 10100 24064
rect 10876 24012 10928 24064
rect 12624 24012 12676 24064
rect 14096 24080 14148 24132
rect 14464 24123 14516 24132
rect 14464 24089 14473 24123
rect 14473 24089 14507 24123
rect 14507 24089 14516 24123
rect 14464 24080 14516 24089
rect 15936 24080 15988 24132
rect 16580 24123 16632 24132
rect 16580 24089 16589 24123
rect 16589 24089 16623 24123
rect 16623 24089 16632 24123
rect 18788 24148 18840 24200
rect 19248 24148 19300 24200
rect 16580 24080 16632 24089
rect 17960 24080 18012 24132
rect 18052 24123 18104 24132
rect 18052 24089 18061 24123
rect 18061 24089 18095 24123
rect 18095 24089 18104 24123
rect 18052 24080 18104 24089
rect 24676 24080 24728 24132
rect 34796 24080 34848 24132
rect 13820 24012 13872 24064
rect 16120 24012 16172 24064
rect 20260 24012 20312 24064
rect 21088 24012 21140 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 2228 23808 2280 23860
rect 3240 23808 3292 23860
rect 5816 23808 5868 23860
rect 6460 23808 6512 23860
rect 7104 23808 7156 23860
rect 6828 23740 6880 23792
rect 10048 23808 10100 23860
rect 8944 23783 8996 23792
rect 8944 23749 8953 23783
rect 8953 23749 8987 23783
rect 8987 23749 8996 23783
rect 8944 23740 8996 23749
rect 9496 23783 9548 23792
rect 9496 23749 9505 23783
rect 9505 23749 9539 23783
rect 9539 23749 9548 23783
rect 11796 23808 11848 23860
rect 10968 23783 11020 23792
rect 9496 23740 9548 23749
rect 10968 23749 10977 23783
rect 10977 23749 11011 23783
rect 11011 23749 11020 23783
rect 10968 23740 11020 23749
rect 11060 23783 11112 23792
rect 11060 23749 11069 23783
rect 11069 23749 11103 23783
rect 11103 23749 11112 23783
rect 13820 23808 13872 23860
rect 14096 23808 14148 23860
rect 27804 23851 27856 23860
rect 27804 23817 27813 23851
rect 27813 23817 27847 23851
rect 27847 23817 27856 23851
rect 27804 23808 27856 23817
rect 11060 23740 11112 23749
rect 12808 23783 12860 23792
rect 12808 23749 12817 23783
rect 12817 23749 12851 23783
rect 12851 23749 12860 23783
rect 12808 23740 12860 23749
rect 2044 23604 2096 23656
rect 3792 23672 3844 23724
rect 7012 23672 7064 23724
rect 5356 23647 5408 23656
rect 1676 23536 1728 23588
rect 5356 23613 5365 23647
rect 5365 23613 5399 23647
rect 5399 23613 5408 23647
rect 5356 23604 5408 23613
rect 5724 23647 5776 23656
rect 5724 23613 5733 23647
rect 5733 23613 5767 23647
rect 5767 23613 5776 23647
rect 5724 23604 5776 23613
rect 8024 23604 8076 23656
rect 3240 23536 3292 23588
rect 3516 23536 3568 23588
rect 4804 23536 4856 23588
rect 8668 23536 8720 23588
rect 8944 23604 8996 23656
rect 10416 23604 10468 23656
rect 11336 23604 11388 23656
rect 11704 23604 11756 23656
rect 12348 23604 12400 23656
rect 12440 23604 12492 23656
rect 15936 23740 15988 23792
rect 16120 23783 16172 23792
rect 16120 23749 16129 23783
rect 16129 23749 16163 23783
rect 16163 23749 16172 23783
rect 16120 23740 16172 23749
rect 17040 23783 17092 23792
rect 17040 23749 17049 23783
rect 17049 23749 17083 23783
rect 17083 23749 17092 23783
rect 17040 23740 17092 23749
rect 17408 23740 17460 23792
rect 20260 23783 20312 23792
rect 20260 23749 20269 23783
rect 20269 23749 20303 23783
rect 20303 23749 20312 23783
rect 20260 23740 20312 23749
rect 13084 23672 13136 23724
rect 18788 23672 18840 23724
rect 27620 23715 27672 23724
rect 14924 23604 14976 23656
rect 16212 23647 16264 23656
rect 10508 23536 10560 23588
rect 11796 23536 11848 23588
rect 16212 23613 16221 23647
rect 16221 23613 16255 23647
rect 16255 23613 16264 23647
rect 16212 23604 16264 23613
rect 17224 23604 17276 23656
rect 19524 23604 19576 23656
rect 21272 23604 21324 23656
rect 3884 23468 3936 23520
rect 5448 23468 5500 23520
rect 14832 23468 14884 23520
rect 17500 23468 17552 23520
rect 19616 23468 19668 23520
rect 27620 23681 27629 23715
rect 27629 23681 27663 23715
rect 27663 23681 27672 23715
rect 27620 23672 27672 23681
rect 23756 23468 23808 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2412 23264 2464 23316
rect 3516 23264 3568 23316
rect 5816 23264 5868 23316
rect 6368 23264 6420 23316
rect 2964 23128 3016 23180
rect 2504 23060 2556 23112
rect 2780 23060 2832 23112
rect 7748 23128 7800 23180
rect 10416 23196 10468 23248
rect 10600 23264 10652 23316
rect 10876 23264 10928 23316
rect 11244 23196 11296 23248
rect 8392 23103 8444 23112
rect 4896 22992 4948 23044
rect 3884 22924 3936 22976
rect 5540 22924 5592 22976
rect 6276 22924 6328 22976
rect 7196 22992 7248 23044
rect 8392 23069 8401 23103
rect 8401 23069 8435 23103
rect 8435 23069 8444 23103
rect 8392 23060 8444 23069
rect 10600 23128 10652 23180
rect 16672 23264 16724 23316
rect 16856 23264 16908 23316
rect 24676 23307 24728 23316
rect 24676 23273 24685 23307
rect 24685 23273 24719 23307
rect 24719 23273 24728 23307
rect 24676 23264 24728 23273
rect 11612 23196 11664 23248
rect 12256 23196 12308 23248
rect 12348 23196 12400 23248
rect 14280 23196 14332 23248
rect 17776 23196 17828 23248
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 13452 23128 13504 23180
rect 15108 23128 15160 23180
rect 16580 23128 16632 23180
rect 19524 23171 19576 23180
rect 19524 23137 19533 23171
rect 19533 23137 19567 23171
rect 19567 23137 19576 23171
rect 19524 23128 19576 23137
rect 14372 23103 14424 23112
rect 8116 22924 8168 22976
rect 9496 22967 9548 22976
rect 9496 22933 9505 22967
rect 9505 22933 9539 22967
rect 9539 22933 9548 22967
rect 9496 22924 9548 22933
rect 9588 22924 9640 22976
rect 11244 22992 11296 23044
rect 11428 22992 11480 23044
rect 11520 23035 11572 23044
rect 11520 23001 11529 23035
rect 11529 23001 11563 23035
rect 11563 23001 11572 23035
rect 11520 22992 11572 23001
rect 12164 22992 12216 23044
rect 14372 23069 14381 23103
rect 14381 23069 14415 23103
rect 14415 23069 14424 23103
rect 14372 23060 14424 23069
rect 14740 23060 14792 23112
rect 13360 22992 13412 23044
rect 13544 23035 13596 23044
rect 13544 23001 13553 23035
rect 13553 23001 13587 23035
rect 13587 23001 13596 23035
rect 13544 22992 13596 23001
rect 16488 23060 16540 23112
rect 17316 23103 17368 23112
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17316 23060 17368 23069
rect 17868 23060 17920 23112
rect 23756 23103 23808 23112
rect 23756 23069 23765 23103
rect 23765 23069 23799 23103
rect 23799 23069 23808 23103
rect 23756 23060 23808 23069
rect 24676 23060 24728 23112
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 19616 23035 19668 23044
rect 19616 23001 19625 23035
rect 19625 23001 19659 23035
rect 19659 23001 19668 23035
rect 19616 22992 19668 23001
rect 18788 22967 18840 22976
rect 18788 22933 18797 22967
rect 18797 22933 18831 22967
rect 18831 22933 18840 22967
rect 18788 22924 18840 22933
rect 23664 22967 23716 22976
rect 23664 22933 23673 22967
rect 23673 22933 23707 22967
rect 23707 22933 23716 22967
rect 23664 22924 23716 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1676 22720 1728 22772
rect 4988 22720 5040 22772
rect 8944 22720 8996 22772
rect 9496 22720 9548 22772
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 2780 22652 2832 22704
rect 6000 22652 6052 22704
rect 6276 22652 6328 22704
rect 7288 22652 7340 22704
rect 8024 22652 8076 22704
rect 9864 22652 9916 22704
rect 11060 22652 11112 22704
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 4896 22584 4948 22593
rect 7472 22584 7524 22636
rect 10232 22584 10284 22636
rect 4896 22448 4948 22500
rect 5264 22448 5316 22500
rect 7104 22516 7156 22568
rect 7196 22516 7248 22568
rect 6552 22448 6604 22500
rect 10324 22516 10376 22568
rect 10600 22584 10652 22636
rect 11980 22584 12032 22636
rect 10876 22516 10928 22568
rect 12256 22652 12308 22704
rect 13360 22652 13412 22704
rect 14464 22652 14516 22704
rect 16212 22720 16264 22772
rect 18052 22720 18104 22772
rect 13728 22627 13780 22636
rect 13728 22593 13737 22627
rect 13737 22593 13771 22627
rect 13771 22593 13780 22627
rect 13728 22584 13780 22593
rect 14924 22559 14976 22568
rect 14924 22525 14933 22559
rect 14933 22525 14967 22559
rect 14967 22525 14976 22559
rect 14924 22516 14976 22525
rect 17960 22516 18012 22568
rect 7380 22380 7432 22432
rect 7932 22380 7984 22432
rect 8300 22380 8352 22432
rect 9036 22380 9088 22432
rect 9772 22448 9824 22500
rect 10600 22448 10652 22500
rect 13176 22448 13228 22500
rect 13360 22448 13412 22500
rect 13728 22448 13780 22500
rect 15108 22448 15160 22500
rect 21180 22652 21232 22704
rect 11060 22423 11112 22432
rect 11060 22389 11069 22423
rect 11069 22389 11103 22423
rect 11103 22389 11112 22423
rect 11060 22380 11112 22389
rect 11152 22380 11204 22432
rect 12348 22380 12400 22432
rect 13084 22380 13136 22432
rect 14924 22380 14976 22432
rect 15476 22380 15528 22432
rect 16764 22380 16816 22432
rect 20260 22584 20312 22636
rect 24860 22584 24912 22636
rect 36268 22491 36320 22500
rect 36268 22457 36277 22491
rect 36277 22457 36311 22491
rect 36311 22457 36320 22491
rect 36268 22448 36320 22457
rect 19616 22423 19668 22432
rect 19616 22389 19625 22423
rect 19625 22389 19659 22423
rect 19659 22389 19668 22423
rect 19616 22380 19668 22389
rect 20260 22423 20312 22432
rect 20260 22389 20269 22423
rect 20269 22389 20303 22423
rect 20303 22389 20312 22423
rect 20260 22380 20312 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 4988 22176 5040 22228
rect 7104 22176 7156 22228
rect 3240 22040 3292 22092
rect 2320 21972 2372 22024
rect 2780 21972 2832 22024
rect 5264 21904 5316 21956
rect 7196 22040 7248 22092
rect 7932 22176 7984 22228
rect 9496 22176 9548 22228
rect 11152 22176 11204 22228
rect 11520 22176 11572 22228
rect 13544 22176 13596 22228
rect 9128 22108 9180 22160
rect 9680 22108 9732 22160
rect 9772 22108 9824 22160
rect 7656 21972 7708 22024
rect 8116 21972 8168 22024
rect 9220 21972 9272 22024
rect 9496 21972 9548 22024
rect 6552 21947 6604 21956
rect 6552 21913 6561 21947
rect 6561 21913 6595 21947
rect 6595 21913 6604 21947
rect 6552 21904 6604 21913
rect 1676 21879 1728 21888
rect 1676 21845 1685 21879
rect 1685 21845 1719 21879
rect 1719 21845 1728 21879
rect 1676 21836 1728 21845
rect 3056 21836 3108 21888
rect 3240 21836 3292 21888
rect 4988 21836 5040 21888
rect 6460 21836 6512 21888
rect 8576 21879 8628 21888
rect 8576 21845 8585 21879
rect 8585 21845 8619 21879
rect 8619 21845 8628 21879
rect 8576 21836 8628 21845
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 9404 21836 9456 21888
rect 9772 21904 9824 21956
rect 10784 22040 10836 22092
rect 10416 21972 10468 22024
rect 11244 21972 11296 22024
rect 13636 22040 13688 22092
rect 13728 22083 13780 22092
rect 13728 22049 13737 22083
rect 13737 22049 13771 22083
rect 13771 22049 13780 22083
rect 14924 22176 14976 22228
rect 15476 22176 15528 22228
rect 19616 22176 19668 22228
rect 13728 22040 13780 22049
rect 10876 21904 10928 21956
rect 11980 21972 12032 22024
rect 14096 21972 14148 22024
rect 18052 22108 18104 22160
rect 18604 22108 18656 22160
rect 14464 22083 14516 22092
rect 14464 22049 14473 22083
rect 14473 22049 14507 22083
rect 14507 22049 14516 22083
rect 14464 22040 14516 22049
rect 14924 22083 14976 22092
rect 14924 22049 14933 22083
rect 14933 22049 14967 22083
rect 14967 22049 14976 22083
rect 14924 22040 14976 22049
rect 15200 22040 15252 22092
rect 15936 22040 15988 22092
rect 16212 21972 16264 22024
rect 20720 21972 20772 22024
rect 35900 21972 35952 22024
rect 15200 21904 15252 21956
rect 17132 21947 17184 21956
rect 17132 21913 17141 21947
rect 17141 21913 17175 21947
rect 17175 21913 17184 21947
rect 17132 21904 17184 21913
rect 17224 21947 17276 21956
rect 17224 21913 17233 21947
rect 17233 21913 17267 21947
rect 17267 21913 17276 21947
rect 17224 21904 17276 21913
rect 18236 21947 18288 21956
rect 18236 21913 18245 21947
rect 18245 21913 18279 21947
rect 18279 21913 18288 21947
rect 18236 21904 18288 21913
rect 10048 21836 10100 21888
rect 12900 21836 12952 21888
rect 15568 21879 15620 21888
rect 15568 21845 15577 21879
rect 15577 21845 15611 21879
rect 15611 21845 15620 21879
rect 15568 21836 15620 21845
rect 17960 21836 18012 21888
rect 19248 21904 19300 21956
rect 22008 21904 22060 21956
rect 20720 21879 20772 21888
rect 20720 21845 20729 21879
rect 20729 21845 20763 21879
rect 20763 21845 20772 21879
rect 20720 21836 20772 21845
rect 21272 21836 21324 21888
rect 21824 21836 21876 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 6828 21675 6880 21684
rect 6828 21641 6837 21675
rect 6837 21641 6871 21675
rect 6871 21641 6880 21675
rect 6828 21632 6880 21641
rect 11888 21632 11940 21684
rect 12624 21675 12676 21684
rect 12624 21641 12633 21675
rect 12633 21641 12667 21675
rect 12667 21641 12676 21675
rect 12624 21632 12676 21641
rect 7564 21607 7616 21616
rect 7564 21573 7573 21607
rect 7573 21573 7607 21607
rect 7607 21573 7616 21607
rect 7564 21564 7616 21573
rect 10416 21564 10468 21616
rect 10692 21564 10744 21616
rect 1860 21539 1912 21548
rect 1860 21505 1869 21539
rect 1869 21505 1903 21539
rect 1903 21505 1912 21539
rect 1860 21496 1912 21505
rect 8944 21496 8996 21548
rect 10600 21496 10652 21548
rect 10876 21496 10928 21548
rect 11152 21564 11204 21616
rect 13636 21564 13688 21616
rect 14188 21564 14240 21616
rect 14464 21607 14516 21616
rect 14464 21573 14473 21607
rect 14473 21573 14507 21607
rect 14507 21573 14516 21607
rect 14464 21564 14516 21573
rect 17040 21632 17092 21684
rect 15108 21607 15160 21616
rect 15108 21573 15117 21607
rect 15117 21573 15151 21607
rect 15151 21573 15160 21607
rect 15108 21564 15160 21573
rect 15384 21564 15436 21616
rect 16120 21607 16172 21616
rect 16120 21573 16129 21607
rect 16129 21573 16163 21607
rect 16163 21573 16172 21607
rect 16120 21564 16172 21573
rect 16212 21564 16264 21616
rect 12532 21496 12584 21548
rect 16856 21539 16908 21548
rect 16856 21505 16865 21539
rect 16865 21505 16899 21539
rect 16899 21505 16908 21539
rect 16856 21496 16908 21505
rect 36268 21539 36320 21548
rect 36268 21505 36277 21539
rect 36277 21505 36311 21539
rect 36311 21505 36320 21539
rect 36268 21496 36320 21505
rect 2780 21428 2832 21480
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 5448 21428 5500 21480
rect 6828 21428 6880 21480
rect 7196 21428 7248 21480
rect 8760 21428 8812 21480
rect 9036 21428 9088 21480
rect 9404 21428 9456 21480
rect 4620 21360 4672 21412
rect 1676 21335 1728 21344
rect 1676 21301 1685 21335
rect 1685 21301 1719 21335
rect 1719 21301 1728 21335
rect 1676 21292 1728 21301
rect 2872 21335 2924 21344
rect 2872 21301 2881 21335
rect 2881 21301 2915 21335
rect 2915 21301 2924 21335
rect 2872 21292 2924 21301
rect 8668 21360 8720 21412
rect 12348 21360 12400 21412
rect 13728 21428 13780 21480
rect 14280 21428 14332 21480
rect 14464 21428 14516 21480
rect 19432 21428 19484 21480
rect 12716 21292 12768 21344
rect 14004 21360 14056 21412
rect 14648 21360 14700 21412
rect 15016 21360 15068 21412
rect 18788 21360 18840 21412
rect 21916 21360 21968 21412
rect 35992 21360 36044 21412
rect 16856 21292 16908 21344
rect 17592 21335 17644 21344
rect 17592 21301 17601 21335
rect 17601 21301 17635 21335
rect 17635 21301 17644 21335
rect 17592 21292 17644 21301
rect 17868 21292 17920 21344
rect 36176 21335 36228 21344
rect 36176 21301 36185 21335
rect 36185 21301 36219 21335
rect 36219 21301 36228 21335
rect 36176 21292 36228 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2780 21088 2832 21140
rect 2872 21088 2924 21140
rect 8392 21088 8444 21140
rect 9128 21088 9180 21140
rect 10968 21131 11020 21140
rect 10968 21097 10977 21131
rect 10977 21097 11011 21131
rect 11011 21097 11020 21131
rect 10968 21088 11020 21097
rect 12256 21131 12308 21140
rect 12256 21097 12265 21131
rect 12265 21097 12299 21131
rect 12299 21097 12308 21131
rect 12256 21088 12308 21097
rect 8760 21020 8812 21072
rect 9404 21020 9456 21072
rect 11152 21020 11204 21072
rect 4988 20952 5040 21004
rect 5080 20952 5132 21004
rect 6460 20952 6512 21004
rect 6828 20952 6880 21004
rect 8944 20952 8996 21004
rect 9496 20952 9548 21004
rect 15016 21088 15068 21140
rect 18236 21088 18288 21140
rect 18788 21088 18840 21140
rect 2780 20884 2832 20936
rect 6552 20927 6604 20936
rect 6552 20893 6561 20927
rect 6561 20893 6595 20927
rect 6595 20893 6604 20927
rect 6552 20884 6604 20893
rect 3424 20859 3476 20868
rect 3424 20825 3433 20859
rect 3433 20825 3467 20859
rect 3467 20825 3476 20859
rect 3424 20816 3476 20825
rect 4252 20816 4304 20868
rect 6000 20816 6052 20868
rect 6460 20816 6512 20868
rect 8208 20816 8260 20868
rect 8668 20816 8720 20868
rect 9956 20884 10008 20936
rect 12440 20952 12492 21004
rect 12992 20952 13044 21004
rect 13360 20952 13412 21004
rect 15384 21020 15436 21072
rect 16212 21020 16264 21072
rect 16488 20952 16540 21004
rect 1860 20748 1912 20800
rect 9404 20816 9456 20868
rect 11244 20884 11296 20936
rect 10968 20816 11020 20868
rect 13636 20884 13688 20936
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 16396 20927 16448 20936
rect 14556 20884 14608 20893
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 16396 20884 16448 20893
rect 16856 20927 16908 20936
rect 16856 20893 16865 20927
rect 16865 20893 16899 20927
rect 16899 20893 16908 20927
rect 16856 20884 16908 20893
rect 13084 20816 13136 20868
rect 8944 20748 8996 20800
rect 11244 20748 11296 20800
rect 11888 20748 11940 20800
rect 12716 20748 12768 20800
rect 15384 20816 15436 20868
rect 15568 20859 15620 20868
rect 15568 20825 15577 20859
rect 15577 20825 15611 20859
rect 15611 20825 15620 20859
rect 15568 20816 15620 20825
rect 19248 20816 19300 20868
rect 16304 20791 16356 20800
rect 16304 20757 16313 20791
rect 16313 20757 16347 20791
rect 16347 20757 16356 20791
rect 16304 20748 16356 20757
rect 19340 20748 19392 20800
rect 21824 20816 21876 20868
rect 36176 20748 36228 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 2780 20544 2832 20596
rect 3424 20587 3476 20596
rect 3424 20553 3433 20587
rect 3433 20553 3467 20587
rect 3467 20553 3476 20587
rect 3424 20544 3476 20553
rect 10232 20544 10284 20596
rect 10416 20587 10468 20596
rect 10416 20553 10425 20587
rect 10425 20553 10459 20587
rect 10459 20553 10468 20587
rect 10416 20544 10468 20553
rect 13728 20544 13780 20596
rect 4252 20519 4304 20528
rect 4252 20485 4261 20519
rect 4261 20485 4295 20519
rect 4295 20485 4304 20519
rect 4252 20476 4304 20485
rect 5356 20476 5408 20528
rect 5540 20476 5592 20528
rect 6460 20476 6512 20528
rect 6828 20519 6880 20528
rect 6828 20485 6837 20519
rect 6837 20485 6871 20519
rect 6871 20485 6880 20519
rect 6828 20476 6880 20485
rect 6920 20476 6972 20528
rect 7472 20476 7524 20528
rect 10784 20476 10836 20528
rect 12440 20476 12492 20528
rect 12900 20519 12952 20528
rect 12900 20485 12909 20519
rect 12909 20485 12943 20519
rect 12943 20485 12952 20519
rect 12900 20476 12952 20485
rect 14924 20544 14976 20596
rect 15200 20587 15252 20596
rect 15200 20553 15209 20587
rect 15209 20553 15243 20587
rect 15243 20553 15252 20587
rect 15200 20544 15252 20553
rect 15660 20544 15712 20596
rect 15108 20476 15160 20528
rect 16764 20476 16816 20528
rect 9128 20408 9180 20460
rect 9772 20408 9824 20460
rect 10048 20408 10100 20460
rect 10324 20408 10376 20460
rect 10600 20408 10652 20460
rect 10692 20408 10744 20460
rect 12348 20408 12400 20460
rect 15292 20451 15344 20460
rect 15292 20417 15301 20451
rect 15301 20417 15335 20451
rect 15335 20417 15344 20451
rect 15292 20408 15344 20417
rect 16580 20408 16632 20460
rect 23296 20544 23348 20596
rect 36084 20544 36136 20596
rect 20260 20408 20312 20460
rect 2964 20340 3016 20392
rect 3332 20340 3384 20392
rect 5908 20383 5960 20392
rect 5908 20349 5917 20383
rect 5917 20349 5951 20383
rect 5951 20349 5960 20383
rect 5908 20340 5960 20349
rect 6552 20340 6604 20392
rect 7196 20340 7248 20392
rect 8760 20340 8812 20392
rect 8852 20340 8904 20392
rect 11796 20340 11848 20392
rect 12532 20340 12584 20392
rect 13452 20340 13504 20392
rect 14280 20272 14332 20324
rect 6736 20204 6788 20256
rect 9404 20204 9456 20256
rect 10048 20204 10100 20256
rect 12624 20204 12676 20256
rect 12716 20204 12768 20256
rect 16028 20315 16080 20324
rect 16028 20281 16037 20315
rect 16037 20281 16071 20315
rect 16071 20281 16080 20315
rect 16028 20272 16080 20281
rect 19616 20272 19668 20324
rect 14924 20204 14976 20256
rect 17224 20204 17276 20256
rect 18420 20204 18472 20256
rect 34520 20204 34572 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 1768 20000 1820 20052
rect 2596 20000 2648 20052
rect 3516 20000 3568 20052
rect 6828 20000 6880 20052
rect 7564 20000 7616 20052
rect 7656 20000 7708 20052
rect 8484 20000 8536 20052
rect 8668 20000 8720 20052
rect 9864 20043 9916 20052
rect 9864 20009 9873 20043
rect 9873 20009 9907 20043
rect 9907 20009 9916 20043
rect 9864 20000 9916 20009
rect 10140 20000 10192 20052
rect 2780 19864 2832 19916
rect 4068 19864 4120 19916
rect 4896 19864 4948 19916
rect 5908 19864 5960 19916
rect 9036 19932 9088 19984
rect 9220 19932 9272 19984
rect 7748 19864 7800 19916
rect 11428 19864 11480 19916
rect 9128 19796 9180 19848
rect 9956 19839 10008 19848
rect 2688 19728 2740 19780
rect 6460 19660 6512 19712
rect 6736 19728 6788 19780
rect 9956 19805 9965 19839
rect 9965 19805 9999 19839
rect 9999 19805 10008 19839
rect 9956 19796 10008 19805
rect 10416 19728 10468 19780
rect 10876 19796 10928 19848
rect 11980 19932 12032 19984
rect 13820 20000 13872 20052
rect 15108 20043 15160 20052
rect 15108 20009 15117 20043
rect 15117 20009 15151 20043
rect 15151 20009 15160 20043
rect 15108 20000 15160 20009
rect 16856 20000 16908 20052
rect 17132 20000 17184 20052
rect 20260 20000 20312 20052
rect 36636 20000 36688 20052
rect 11796 19907 11848 19916
rect 11796 19873 11805 19907
rect 11805 19873 11839 19907
rect 11839 19873 11848 19907
rect 11796 19864 11848 19873
rect 12164 19864 12216 19916
rect 13452 19864 13504 19916
rect 14280 19864 14332 19916
rect 14464 19839 14516 19848
rect 8300 19660 8352 19712
rect 9036 19660 9088 19712
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 11888 19771 11940 19780
rect 11888 19737 11897 19771
rect 11897 19737 11931 19771
rect 11931 19737 11940 19771
rect 11888 19728 11940 19737
rect 12072 19728 12124 19780
rect 13452 19771 13504 19780
rect 13084 19660 13136 19712
rect 13452 19737 13461 19771
rect 13461 19737 13495 19771
rect 13495 19737 13504 19771
rect 13452 19728 13504 19737
rect 13728 19728 13780 19780
rect 17316 19932 17368 19984
rect 19064 19932 19116 19984
rect 19432 19932 19484 19984
rect 20444 19864 20496 19916
rect 14372 19660 14424 19712
rect 15200 19660 15252 19712
rect 18420 19796 18472 19848
rect 22468 19839 22520 19848
rect 22468 19805 22477 19839
rect 22477 19805 22511 19839
rect 22511 19805 22520 19839
rect 22928 19839 22980 19848
rect 22468 19796 22520 19805
rect 22928 19805 22937 19839
rect 22937 19805 22971 19839
rect 22971 19805 22980 19839
rect 22928 19796 22980 19805
rect 18604 19728 18656 19780
rect 19616 19771 19668 19780
rect 19616 19737 19625 19771
rect 19625 19737 19659 19771
rect 19659 19737 19668 19771
rect 20168 19771 20220 19780
rect 19616 19728 19668 19737
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 20536 19728 20588 19780
rect 16580 19660 16632 19712
rect 18144 19703 18196 19712
rect 18144 19669 18153 19703
rect 18153 19669 18187 19703
rect 18187 19669 18196 19703
rect 18144 19660 18196 19669
rect 22192 19660 22244 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3516 19388 3568 19440
rect 5540 19456 5592 19508
rect 5816 19456 5868 19508
rect 6460 19456 6512 19508
rect 7656 19456 7708 19508
rect 7472 19388 7524 19440
rect 8576 19456 8628 19508
rect 8760 19456 8812 19508
rect 9588 19388 9640 19440
rect 12624 19431 12676 19440
rect 1584 19363 1636 19372
rect 1584 19329 1593 19363
rect 1593 19329 1627 19363
rect 1627 19329 1636 19363
rect 1584 19320 1636 19329
rect 4068 19320 4120 19372
rect 6920 19363 6972 19372
rect 6920 19329 6929 19363
rect 6929 19329 6963 19363
rect 6963 19329 6972 19363
rect 6920 19320 6972 19329
rect 7104 19320 7156 19372
rect 9404 19320 9456 19372
rect 10416 19320 10468 19372
rect 1952 19252 2004 19304
rect 4528 19295 4580 19304
rect 4528 19261 4537 19295
rect 4537 19261 4571 19295
rect 4571 19261 4580 19295
rect 4528 19252 4580 19261
rect 5264 19252 5316 19304
rect 7196 19252 7248 19304
rect 7288 19252 7340 19304
rect 11428 19320 11480 19372
rect 12072 19320 12124 19372
rect 5540 19184 5592 19236
rect 7012 19184 7064 19236
rect 7104 19184 7156 19236
rect 7380 19184 7432 19236
rect 8760 19184 8812 19236
rect 11888 19184 11940 19236
rect 12624 19397 12633 19431
rect 12633 19397 12667 19431
rect 12667 19397 12676 19431
rect 12624 19388 12676 19397
rect 13452 19456 13504 19508
rect 16120 19456 16172 19508
rect 14832 19388 14884 19440
rect 13544 19320 13596 19372
rect 14648 19320 14700 19372
rect 18144 19388 18196 19440
rect 19340 19456 19392 19508
rect 18788 19388 18840 19440
rect 21272 19388 21324 19440
rect 22192 19431 22244 19440
rect 22192 19397 22201 19431
rect 22201 19397 22235 19431
rect 22235 19397 22244 19431
rect 22192 19388 22244 19397
rect 15016 19363 15068 19372
rect 15016 19329 15025 19363
rect 15025 19329 15059 19363
rect 15059 19329 15068 19363
rect 15016 19320 15068 19329
rect 15936 19320 15988 19372
rect 16120 19320 16172 19372
rect 16396 19320 16448 19372
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 19064 19363 19116 19372
rect 19064 19329 19073 19363
rect 19073 19329 19107 19363
rect 19107 19329 19116 19363
rect 19064 19320 19116 19329
rect 19708 19320 19760 19372
rect 35900 19363 35952 19372
rect 35900 19329 35909 19363
rect 35909 19329 35943 19363
rect 35943 19329 35952 19363
rect 35900 19320 35952 19329
rect 12716 19252 12768 19304
rect 14004 19252 14056 19304
rect 14740 19252 14792 19304
rect 14924 19252 14976 19304
rect 16948 19295 17000 19304
rect 12440 19184 12492 19236
rect 12808 19184 12860 19236
rect 16120 19184 16172 19236
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 19984 19252 20036 19304
rect 21088 19295 21140 19304
rect 21088 19261 21097 19295
rect 21097 19261 21131 19295
rect 21131 19261 21140 19295
rect 21088 19252 21140 19261
rect 22100 19295 22152 19304
rect 22100 19261 22109 19295
rect 22109 19261 22143 19295
rect 22143 19261 22152 19295
rect 22100 19252 22152 19261
rect 2504 19116 2556 19168
rect 4896 19116 4948 19168
rect 5264 19116 5316 19168
rect 9312 19116 9364 19168
rect 10416 19159 10468 19168
rect 10416 19125 10425 19159
rect 10425 19125 10459 19159
rect 10459 19125 10468 19159
rect 10416 19116 10468 19125
rect 12072 19116 12124 19168
rect 15384 19116 15436 19168
rect 15844 19116 15896 19168
rect 36084 19159 36136 19168
rect 36084 19125 36093 19159
rect 36093 19125 36127 19159
rect 36127 19125 36136 19159
rect 36084 19116 36136 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1400 18912 1452 18964
rect 6092 18912 6144 18964
rect 7012 18912 7064 18964
rect 7196 18912 7248 18964
rect 14372 18955 14424 18964
rect 14372 18921 14381 18955
rect 14381 18921 14415 18955
rect 14415 18921 14424 18955
rect 14372 18912 14424 18921
rect 15292 18912 15344 18964
rect 16580 18912 16632 18964
rect 29828 18912 29880 18964
rect 4068 18776 4120 18828
rect 5172 18776 5224 18828
rect 5632 18776 5684 18828
rect 6368 18844 6420 18896
rect 7288 18776 7340 18828
rect 9864 18776 9916 18828
rect 13544 18844 13596 18896
rect 14096 18844 14148 18896
rect 9588 18751 9640 18760
rect 9588 18717 9597 18751
rect 9597 18717 9631 18751
rect 9631 18717 9640 18751
rect 9588 18708 9640 18717
rect 9956 18708 10008 18760
rect 10600 18708 10652 18760
rect 11796 18776 11848 18828
rect 15200 18776 15252 18828
rect 15476 18819 15528 18828
rect 15476 18785 15485 18819
rect 15485 18785 15519 18819
rect 15519 18785 15528 18819
rect 15476 18776 15528 18785
rect 14280 18708 14332 18760
rect 16488 18844 16540 18896
rect 16948 18776 17000 18828
rect 20628 18844 20680 18896
rect 24860 18844 24912 18896
rect 20168 18776 20220 18828
rect 21824 18819 21876 18828
rect 21824 18785 21833 18819
rect 21833 18785 21867 18819
rect 21867 18785 21876 18819
rect 21824 18776 21876 18785
rect 5264 18640 5316 18692
rect 7840 18640 7892 18692
rect 8300 18683 8352 18692
rect 8300 18649 8309 18683
rect 8309 18649 8343 18683
rect 8343 18649 8352 18683
rect 8300 18640 8352 18649
rect 10416 18640 10468 18692
rect 10140 18615 10192 18624
rect 10140 18581 10149 18615
rect 10149 18581 10183 18615
rect 10183 18581 10192 18615
rect 10140 18572 10192 18581
rect 12164 18640 12216 18692
rect 13084 18683 13136 18692
rect 13084 18649 13093 18683
rect 13093 18649 13127 18683
rect 13127 18649 13136 18683
rect 13084 18640 13136 18649
rect 14004 18640 14056 18692
rect 15384 18683 15436 18692
rect 15384 18649 15393 18683
rect 15393 18649 15427 18683
rect 15427 18649 15436 18683
rect 15384 18640 15436 18649
rect 17960 18640 18012 18692
rect 18696 18683 18748 18692
rect 18696 18649 18705 18683
rect 18705 18649 18739 18683
rect 18739 18649 18748 18683
rect 18696 18640 18748 18649
rect 18788 18683 18840 18692
rect 18788 18649 18797 18683
rect 18797 18649 18831 18683
rect 18831 18649 18840 18683
rect 18788 18640 18840 18649
rect 18972 18640 19024 18692
rect 12624 18572 12676 18624
rect 15292 18572 15344 18624
rect 20628 18640 20680 18692
rect 21180 18683 21232 18692
rect 21180 18649 21189 18683
rect 21189 18649 21223 18683
rect 21223 18649 21232 18683
rect 21180 18640 21232 18649
rect 19800 18572 19852 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2504 18368 2556 18420
rect 3424 18368 3476 18420
rect 5540 18368 5592 18420
rect 6000 18368 6052 18420
rect 4344 18300 4396 18352
rect 10140 18368 10192 18420
rect 7564 18300 7616 18352
rect 9772 18300 9824 18352
rect 5908 18275 5960 18284
rect 5908 18241 5917 18275
rect 5917 18241 5951 18275
rect 5951 18241 5960 18275
rect 5908 18232 5960 18241
rect 7012 18232 7064 18284
rect 8852 18232 8904 18284
rect 9864 18232 9916 18284
rect 1952 18164 2004 18216
rect 3424 18207 3476 18216
rect 3424 18173 3433 18207
rect 3433 18173 3467 18207
rect 3467 18173 3476 18207
rect 3424 18164 3476 18173
rect 5632 18207 5684 18216
rect 5632 18173 5641 18207
rect 5641 18173 5675 18207
rect 5675 18173 5684 18207
rect 5632 18164 5684 18173
rect 7196 18207 7248 18216
rect 7196 18173 7205 18207
rect 7205 18173 7239 18207
rect 7239 18173 7248 18207
rect 7196 18164 7248 18173
rect 8760 18164 8812 18216
rect 9312 18164 9364 18216
rect 14372 18368 14424 18420
rect 18788 18368 18840 18420
rect 21272 18411 21324 18420
rect 12072 18343 12124 18352
rect 12072 18309 12081 18343
rect 12081 18309 12115 18343
rect 12115 18309 12124 18343
rect 12072 18300 12124 18309
rect 12624 18343 12676 18352
rect 12624 18309 12633 18343
rect 12633 18309 12667 18343
rect 12667 18309 12676 18343
rect 12624 18300 12676 18309
rect 13728 18343 13780 18352
rect 13728 18309 13737 18343
rect 13737 18309 13771 18343
rect 13771 18309 13780 18343
rect 13728 18300 13780 18309
rect 15200 18343 15252 18352
rect 15200 18309 15209 18343
rect 15209 18309 15243 18343
rect 15243 18309 15252 18343
rect 15200 18300 15252 18309
rect 10416 18232 10468 18284
rect 10876 18232 10928 18284
rect 12440 18164 12492 18216
rect 8668 18096 8720 18148
rect 16764 18232 16816 18284
rect 19064 18232 19116 18284
rect 19432 18300 19484 18352
rect 21272 18377 21281 18411
rect 21281 18377 21315 18411
rect 21315 18377 21324 18411
rect 21272 18368 21324 18377
rect 22928 18411 22980 18420
rect 22928 18377 22937 18411
rect 22937 18377 22971 18411
rect 22971 18377 22980 18411
rect 22928 18368 22980 18377
rect 27620 18300 27672 18352
rect 21088 18232 21140 18284
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 22928 18232 22980 18284
rect 34520 18232 34572 18284
rect 36084 18275 36136 18284
rect 36084 18241 36093 18275
rect 36093 18241 36127 18275
rect 36127 18241 36136 18275
rect 36084 18232 36136 18241
rect 13176 18164 13228 18216
rect 13636 18207 13688 18216
rect 13636 18173 13645 18207
rect 13645 18173 13679 18207
rect 13679 18173 13688 18207
rect 13636 18164 13688 18173
rect 15292 18164 15344 18216
rect 19248 18164 19300 18216
rect 20168 18207 20220 18216
rect 20168 18173 20177 18207
rect 20177 18173 20211 18207
rect 20211 18173 20220 18207
rect 20168 18164 20220 18173
rect 20628 18207 20680 18216
rect 20628 18173 20637 18207
rect 20637 18173 20671 18207
rect 20671 18173 20680 18207
rect 20628 18164 20680 18173
rect 21732 18096 21784 18148
rect 6184 18028 6236 18080
rect 11980 18028 12032 18080
rect 17960 18028 18012 18080
rect 19340 18028 19392 18080
rect 19984 18028 20036 18080
rect 22376 18071 22428 18080
rect 22376 18037 22385 18071
rect 22385 18037 22419 18071
rect 22419 18037 22428 18071
rect 22376 18028 22428 18037
rect 36268 18071 36320 18080
rect 36268 18037 36277 18071
rect 36277 18037 36311 18071
rect 36311 18037 36320 18071
rect 36268 18028 36320 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 8484 17867 8536 17876
rect 3516 17756 3568 17808
rect 8484 17833 8493 17867
rect 8493 17833 8527 17867
rect 8527 17833 8536 17867
rect 8484 17824 8536 17833
rect 10784 17867 10836 17876
rect 10784 17833 10793 17867
rect 10793 17833 10827 17867
rect 10827 17833 10836 17867
rect 10784 17824 10836 17833
rect 12532 17824 12584 17876
rect 2412 17688 2464 17740
rect 4068 17688 4120 17740
rect 4436 17731 4488 17740
rect 4436 17697 4445 17731
rect 4445 17697 4479 17731
rect 4479 17697 4488 17731
rect 4436 17688 4488 17697
rect 6736 17756 6788 17808
rect 8116 17756 8168 17808
rect 10876 17756 10928 17808
rect 19432 17824 19484 17876
rect 22100 17824 22152 17876
rect 6368 17688 6420 17740
rect 6460 17688 6512 17740
rect 7748 17688 7800 17740
rect 10508 17688 10560 17740
rect 12164 17688 12216 17740
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 4712 17595 4764 17604
rect 4712 17561 4721 17595
rect 4721 17561 4755 17595
rect 4755 17561 4764 17595
rect 4712 17552 4764 17561
rect 4804 17484 4856 17536
rect 6644 17552 6696 17604
rect 8852 17620 8904 17672
rect 9588 17663 9640 17672
rect 9588 17629 9597 17663
rect 9597 17629 9631 17663
rect 9631 17629 9640 17663
rect 9588 17620 9640 17629
rect 10416 17620 10468 17672
rect 10600 17620 10652 17672
rect 13268 17688 13320 17740
rect 15200 17688 15252 17740
rect 12716 17620 12768 17672
rect 16764 17756 16816 17808
rect 20168 17756 20220 17808
rect 16396 17688 16448 17740
rect 20536 17731 20588 17740
rect 7288 17552 7340 17604
rect 9680 17552 9732 17604
rect 11612 17595 11664 17604
rect 11612 17561 11621 17595
rect 11621 17561 11655 17595
rect 11655 17561 11664 17595
rect 11612 17552 11664 17561
rect 12624 17552 12676 17604
rect 13084 17595 13136 17604
rect 13084 17561 13093 17595
rect 13093 17561 13127 17595
rect 13127 17561 13136 17595
rect 13084 17552 13136 17561
rect 14832 17595 14884 17604
rect 5724 17484 5776 17536
rect 7656 17484 7708 17536
rect 10048 17484 10100 17536
rect 12440 17484 12492 17536
rect 14832 17561 14841 17595
rect 14841 17561 14875 17595
rect 14875 17561 14884 17595
rect 14832 17552 14884 17561
rect 20536 17697 20545 17731
rect 20545 17697 20579 17731
rect 20579 17697 20588 17731
rect 20536 17688 20588 17697
rect 19432 17620 19484 17672
rect 18236 17552 18288 17604
rect 20996 17552 21048 17604
rect 15936 17484 15988 17536
rect 19064 17484 19116 17536
rect 20168 17484 20220 17536
rect 22376 17756 22428 17808
rect 21640 17688 21692 17740
rect 21824 17663 21876 17672
rect 21824 17629 21833 17663
rect 21833 17629 21867 17663
rect 21867 17629 21876 17663
rect 21824 17620 21876 17629
rect 36544 17484 36596 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 3976 17280 4028 17332
rect 1584 17212 1636 17264
rect 1492 17144 1544 17196
rect 2412 17051 2464 17060
rect 2412 17017 2421 17051
rect 2421 17017 2455 17051
rect 2455 17017 2464 17051
rect 2412 17008 2464 17017
rect 3792 17212 3844 17264
rect 5540 17280 5592 17332
rect 6644 17280 6696 17332
rect 7104 17212 7156 17264
rect 7840 17212 7892 17264
rect 9220 17212 9272 17264
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6276 17144 6328 17196
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 2964 17008 3016 17060
rect 3700 17076 3752 17128
rect 3976 17076 4028 17128
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 7288 17076 7340 17085
rect 10232 17280 10284 17332
rect 10416 17280 10468 17332
rect 11612 17280 11664 17332
rect 21640 17280 21692 17332
rect 11888 17255 11940 17264
rect 11888 17221 11897 17255
rect 11897 17221 11931 17255
rect 11931 17221 11940 17255
rect 11888 17212 11940 17221
rect 11980 17212 12032 17264
rect 13636 17212 13688 17264
rect 15384 17255 15436 17264
rect 15384 17221 15393 17255
rect 15393 17221 15427 17255
rect 15427 17221 15436 17255
rect 15384 17212 15436 17221
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 11152 17144 11204 17196
rect 16396 17212 16448 17264
rect 17500 17212 17552 17264
rect 20996 17255 21048 17264
rect 20996 17221 21005 17255
rect 21005 17221 21039 17255
rect 21039 17221 21048 17255
rect 20996 17212 21048 17221
rect 21088 17212 21140 17264
rect 12164 17076 12216 17128
rect 12992 17119 13044 17128
rect 12992 17085 13001 17119
rect 13001 17085 13035 17119
rect 13035 17085 13044 17119
rect 12992 17076 13044 17085
rect 14096 17076 14148 17128
rect 4436 16940 4488 16992
rect 4712 16940 4764 16992
rect 5540 16940 5592 16992
rect 7380 16940 7432 16992
rect 10692 16940 10744 16992
rect 13268 17008 13320 17060
rect 15108 17076 15160 17128
rect 14280 16983 14332 16992
rect 14280 16949 14289 16983
rect 14289 16949 14323 16983
rect 14323 16949 14332 16983
rect 14280 16940 14332 16949
rect 15016 16940 15068 16992
rect 19616 17076 19668 17128
rect 16396 17008 16448 17060
rect 18420 17008 18472 17060
rect 18880 17051 18932 17060
rect 18880 17017 18889 17051
rect 18889 17017 18923 17051
rect 18923 17017 18932 17051
rect 18880 17008 18932 17017
rect 21732 17076 21784 17128
rect 21456 17008 21508 17060
rect 15844 16940 15896 16992
rect 18328 16983 18380 16992
rect 18328 16949 18337 16983
rect 18337 16949 18371 16983
rect 18371 16949 18380 16983
rect 18328 16940 18380 16949
rect 19432 16940 19484 16992
rect 19708 16983 19760 16992
rect 19708 16949 19717 16983
rect 19717 16949 19751 16983
rect 19751 16949 19760 16983
rect 19708 16940 19760 16949
rect 19800 16940 19852 16992
rect 21548 16940 21600 16992
rect 22468 16940 22520 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1676 16736 1728 16788
rect 1860 16736 1912 16788
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 4068 16736 4120 16788
rect 7380 16668 7432 16720
rect 7748 16668 7800 16720
rect 12532 16736 12584 16788
rect 18972 16736 19024 16788
rect 19800 16736 19852 16788
rect 20996 16736 21048 16788
rect 21456 16779 21508 16788
rect 21456 16745 21465 16779
rect 21465 16745 21499 16779
rect 21499 16745 21508 16779
rect 21456 16736 21508 16745
rect 21548 16736 21600 16788
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 3148 16600 3200 16652
rect 3976 16600 4028 16652
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 4252 16600 4304 16609
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 7012 16532 7064 16584
rect 7932 16575 7984 16584
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 8208 16532 8260 16584
rect 8852 16532 8904 16584
rect 18052 16668 18104 16720
rect 19708 16668 19760 16720
rect 20352 16668 20404 16720
rect 21916 16711 21968 16720
rect 12532 16600 12584 16652
rect 13176 16643 13228 16652
rect 13176 16609 13185 16643
rect 13185 16609 13219 16643
rect 13219 16609 13228 16643
rect 13176 16600 13228 16609
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 18328 16600 18380 16652
rect 19616 16600 19668 16652
rect 4896 16464 4948 16516
rect 5080 16464 5132 16516
rect 5724 16464 5776 16516
rect 4528 16396 4580 16448
rect 5172 16396 5224 16448
rect 5356 16396 5408 16448
rect 14648 16532 14700 16584
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 18512 16532 18564 16584
rect 20536 16532 20588 16584
rect 21916 16677 21925 16711
rect 21925 16677 21959 16711
rect 21959 16677 21968 16711
rect 21916 16668 21968 16677
rect 36452 16668 36504 16720
rect 7380 16396 7432 16448
rect 10784 16396 10836 16448
rect 11244 16396 11296 16448
rect 14280 16464 14332 16516
rect 15844 16507 15896 16516
rect 14648 16439 14700 16448
rect 14648 16405 14657 16439
rect 14657 16405 14691 16439
rect 14691 16405 14700 16439
rect 15844 16473 15853 16507
rect 15853 16473 15887 16507
rect 15887 16473 15896 16507
rect 15844 16464 15896 16473
rect 16948 16507 17000 16516
rect 16948 16473 16957 16507
rect 16957 16473 16991 16507
rect 16991 16473 17000 16507
rect 16948 16464 17000 16473
rect 14648 16396 14700 16405
rect 19340 16396 19392 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4896 16192 4948 16244
rect 6920 16192 6972 16244
rect 3240 16124 3292 16176
rect 2688 16056 2740 16108
rect 4988 16056 5040 16108
rect 6736 16124 6788 16176
rect 9036 16192 9088 16244
rect 7380 16124 7432 16176
rect 7656 16167 7708 16176
rect 7656 16133 7665 16167
rect 7665 16133 7699 16167
rect 7699 16133 7708 16167
rect 7656 16124 7708 16133
rect 9312 16124 9364 16176
rect 10232 16124 10284 16176
rect 10692 16124 10744 16176
rect 13728 16192 13780 16244
rect 15384 16192 15436 16244
rect 16948 16235 17000 16244
rect 16948 16201 16957 16235
rect 16957 16201 16991 16235
rect 16991 16201 17000 16235
rect 16948 16192 17000 16201
rect 17224 16192 17276 16244
rect 19892 16192 19944 16244
rect 20536 16192 20588 16244
rect 5540 16056 5592 16108
rect 5724 16056 5776 16108
rect 7012 16056 7064 16108
rect 4528 15988 4580 16040
rect 5172 15988 5224 16040
rect 10784 16056 10836 16108
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 14372 16124 14424 16176
rect 17316 16124 17368 16176
rect 19340 16124 19392 16176
rect 19800 16124 19852 16176
rect 16120 16099 16172 16108
rect 2780 15920 2832 15972
rect 5264 15920 5316 15972
rect 7012 15920 7064 15972
rect 7288 15920 7340 15972
rect 10324 15963 10376 15972
rect 2320 15895 2372 15904
rect 2320 15861 2329 15895
rect 2329 15861 2363 15895
rect 2363 15861 2372 15895
rect 2320 15852 2372 15861
rect 2504 15852 2556 15904
rect 10324 15929 10333 15963
rect 10333 15929 10367 15963
rect 10367 15929 10376 15963
rect 10324 15920 10376 15929
rect 12808 15852 12860 15904
rect 16120 16065 16129 16099
rect 16129 16065 16163 16099
rect 16163 16065 16172 16099
rect 16120 16056 16172 16065
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 22560 16099 22612 16108
rect 22560 16065 22569 16099
rect 22569 16065 22603 16099
rect 22603 16065 22612 16099
rect 22560 16056 22612 16065
rect 36360 16099 36412 16108
rect 12992 15988 13044 16040
rect 14096 15988 14148 16040
rect 14924 15988 14976 16040
rect 15292 16031 15344 16040
rect 15292 15997 15301 16031
rect 15301 15997 15335 16031
rect 15335 15997 15344 16031
rect 15292 15988 15344 15997
rect 16212 15988 16264 16040
rect 16580 15920 16632 15972
rect 20076 15988 20128 16040
rect 20628 15988 20680 16040
rect 20168 15920 20220 15972
rect 16028 15852 16080 15904
rect 17500 15852 17552 15904
rect 18512 15852 18564 15904
rect 18788 15852 18840 15904
rect 36360 16065 36369 16099
rect 36369 16065 36403 16099
rect 36403 16065 36412 16099
rect 36360 16056 36412 16065
rect 35900 15852 35952 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 6460 15648 6512 15700
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 8576 15648 8628 15700
rect 8944 15648 8996 15700
rect 10876 15691 10928 15700
rect 10876 15657 10885 15691
rect 10885 15657 10919 15691
rect 10919 15657 10928 15691
rect 10876 15648 10928 15657
rect 8668 15512 8720 15564
rect 14464 15648 14516 15700
rect 17316 15691 17368 15700
rect 17316 15657 17325 15691
rect 17325 15657 17359 15691
rect 17359 15657 17368 15691
rect 17316 15648 17368 15657
rect 18696 15691 18748 15700
rect 18696 15657 18705 15691
rect 18705 15657 18739 15691
rect 18739 15657 18748 15691
rect 18696 15648 18748 15657
rect 22560 15648 22612 15700
rect 30564 15648 30616 15700
rect 14188 15512 14240 15564
rect 4160 15444 4212 15496
rect 6368 15444 6420 15496
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 10508 15444 10560 15496
rect 14096 15444 14148 15496
rect 19892 15580 19944 15632
rect 20628 15580 20680 15632
rect 15568 15512 15620 15564
rect 16304 15512 16356 15564
rect 20260 15512 20312 15564
rect 1400 15376 1452 15428
rect 6092 15376 6144 15428
rect 4712 15308 4764 15360
rect 4896 15308 4948 15360
rect 7380 15308 7432 15360
rect 9496 15376 9548 15428
rect 11060 15376 11112 15428
rect 10048 15308 10100 15360
rect 12164 15308 12216 15360
rect 12808 15376 12860 15428
rect 13084 15419 13136 15428
rect 13084 15385 13093 15419
rect 13093 15385 13127 15419
rect 13127 15385 13136 15419
rect 13084 15376 13136 15385
rect 12992 15308 13044 15360
rect 15292 15376 15344 15428
rect 15752 15376 15804 15428
rect 17316 15444 17368 15496
rect 18144 15444 18196 15496
rect 17592 15376 17644 15428
rect 18972 15444 19024 15496
rect 19800 15444 19852 15496
rect 20904 15444 20956 15496
rect 16764 15351 16816 15360
rect 16764 15317 16773 15351
rect 16773 15317 16807 15351
rect 16807 15317 16816 15351
rect 16764 15308 16816 15317
rect 17776 15308 17828 15360
rect 18788 15376 18840 15428
rect 20444 15419 20496 15428
rect 20444 15385 20453 15419
rect 20453 15385 20487 15419
rect 20487 15385 20496 15419
rect 20444 15376 20496 15385
rect 22192 15419 22244 15428
rect 22192 15385 22201 15419
rect 22201 15385 22235 15419
rect 22235 15385 22244 15419
rect 22192 15376 22244 15385
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 3056 15104 3108 15156
rect 5356 15104 5408 15156
rect 2872 15036 2924 15088
rect 3424 15036 3476 15088
rect 3792 15036 3844 15088
rect 4068 14968 4120 15020
rect 10324 15104 10376 15156
rect 11060 15104 11112 15156
rect 11888 15104 11940 15156
rect 13268 15104 13320 15156
rect 13452 15104 13504 15156
rect 10968 15079 11020 15088
rect 10968 15045 10977 15079
rect 10977 15045 11011 15079
rect 11011 15045 11020 15079
rect 10968 15036 11020 15045
rect 11336 15036 11388 15088
rect 13636 15036 13688 15088
rect 15108 15104 15160 15156
rect 10416 14968 10468 15020
rect 11244 14968 11296 15020
rect 3976 14900 4028 14952
rect 4160 14900 4212 14952
rect 6920 14900 6972 14952
rect 3884 14832 3936 14884
rect 8300 14900 8352 14952
rect 9404 14900 9456 14952
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 11336 14900 11388 14952
rect 11796 14968 11848 15020
rect 12532 14832 12584 14884
rect 13268 14832 13320 14884
rect 15016 15036 15068 15088
rect 17868 15104 17920 15156
rect 20444 15104 20496 15156
rect 15384 15079 15436 15088
rect 15384 15045 15393 15079
rect 15393 15045 15427 15079
rect 15427 15045 15436 15079
rect 15384 15036 15436 15045
rect 16764 15036 16816 15088
rect 17960 15036 18012 15088
rect 18604 15036 18656 15088
rect 17592 14968 17644 15020
rect 18328 14968 18380 15020
rect 20260 15036 20312 15088
rect 21180 15036 21232 15088
rect 20720 14968 20772 15020
rect 21272 14968 21324 15020
rect 14188 14900 14240 14952
rect 14464 14900 14516 14952
rect 15660 14943 15712 14952
rect 15660 14909 15669 14943
rect 15669 14909 15703 14943
rect 15703 14909 15712 14943
rect 15660 14900 15712 14909
rect 17224 14943 17276 14952
rect 17224 14909 17233 14943
rect 17233 14909 17267 14943
rect 17267 14909 17276 14943
rect 17224 14900 17276 14909
rect 20076 14900 20128 14952
rect 20628 14900 20680 14952
rect 13820 14832 13872 14884
rect 2596 14764 2648 14816
rect 11796 14764 11848 14816
rect 21272 14764 21324 14816
rect 23480 14764 23532 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3608 14560 3660 14612
rect 7012 14560 7064 14612
rect 2964 14492 3016 14544
rect 5724 14492 5776 14544
rect 6184 14492 6236 14544
rect 9404 14560 9456 14612
rect 12532 14560 12584 14612
rect 12992 14603 13044 14612
rect 12992 14569 13001 14603
rect 13001 14569 13035 14603
rect 13035 14569 13044 14603
rect 12992 14560 13044 14569
rect 13636 14603 13688 14612
rect 13636 14569 13645 14603
rect 13645 14569 13679 14603
rect 13679 14569 13688 14603
rect 13636 14560 13688 14569
rect 15016 14603 15068 14612
rect 15016 14569 15025 14603
rect 15025 14569 15059 14603
rect 15059 14569 15068 14603
rect 15016 14560 15068 14569
rect 15292 14560 15344 14612
rect 16120 14560 16172 14612
rect 18788 14603 18840 14612
rect 18788 14569 18797 14603
rect 18797 14569 18831 14603
rect 18831 14569 18840 14603
rect 18788 14560 18840 14569
rect 1584 14424 1636 14476
rect 2044 14424 2096 14476
rect 2412 14424 2464 14476
rect 6828 14424 6880 14476
rect 6920 14424 6972 14476
rect 8576 14467 8628 14476
rect 8576 14433 8585 14467
rect 8585 14433 8619 14467
rect 8619 14433 8628 14467
rect 8576 14424 8628 14433
rect 12348 14424 12400 14476
rect 18052 14467 18104 14476
rect 5356 14356 5408 14408
rect 10784 14356 10836 14408
rect 5264 14288 5316 14340
rect 7012 14288 7064 14340
rect 7840 14288 7892 14340
rect 8300 14331 8352 14340
rect 8300 14297 8309 14331
rect 8309 14297 8343 14331
rect 8343 14297 8352 14331
rect 8300 14288 8352 14297
rect 8760 14288 8812 14340
rect 13360 14356 13412 14408
rect 13544 14356 13596 14408
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14464 14356 14516 14365
rect 18052 14433 18061 14467
rect 18061 14433 18095 14467
rect 18095 14433 18104 14467
rect 18052 14424 18104 14433
rect 19984 14467 20036 14476
rect 19984 14433 19993 14467
rect 19993 14433 20027 14467
rect 20027 14433 20036 14467
rect 19984 14424 20036 14433
rect 22192 14492 22244 14544
rect 20628 14424 20680 14476
rect 3516 14220 3568 14272
rect 4528 14220 4580 14272
rect 5816 14220 5868 14272
rect 11980 14331 12032 14340
rect 11980 14297 11989 14331
rect 11989 14297 12023 14331
rect 12023 14297 12032 14331
rect 11980 14288 12032 14297
rect 12072 14331 12124 14340
rect 12072 14297 12081 14331
rect 12081 14297 12115 14331
rect 12115 14297 12124 14331
rect 16396 14356 16448 14408
rect 12072 14288 12124 14297
rect 9588 14220 9640 14272
rect 10140 14220 10192 14272
rect 10784 14220 10836 14272
rect 13636 14220 13688 14272
rect 15292 14220 15344 14272
rect 20076 14331 20128 14340
rect 20076 14297 20085 14331
rect 20085 14297 20119 14331
rect 20119 14297 20128 14331
rect 20076 14288 20128 14297
rect 21088 14331 21140 14340
rect 17868 14220 17920 14272
rect 21088 14297 21097 14331
rect 21097 14297 21131 14331
rect 21131 14297 21140 14331
rect 21088 14288 21140 14297
rect 21640 14331 21692 14340
rect 21640 14297 21649 14331
rect 21649 14297 21683 14331
rect 21683 14297 21692 14331
rect 21640 14288 21692 14297
rect 21732 14331 21784 14340
rect 21732 14297 21741 14331
rect 21741 14297 21775 14331
rect 21775 14297 21784 14331
rect 21732 14288 21784 14297
rect 22468 14331 22520 14340
rect 22468 14297 22477 14331
rect 22477 14297 22511 14331
rect 22511 14297 22520 14331
rect 22468 14288 22520 14297
rect 22744 14220 22796 14272
rect 35532 14263 35584 14272
rect 35532 14229 35541 14263
rect 35541 14229 35575 14263
rect 35575 14229 35584 14263
rect 36268 14263 36320 14272
rect 35532 14220 35584 14229
rect 36268 14229 36277 14263
rect 36277 14229 36311 14263
rect 36311 14229 36320 14263
rect 36268 14220 36320 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 3976 14016 4028 14068
rect 1860 13948 1912 14000
rect 5172 14016 5224 14068
rect 6828 14016 6880 14068
rect 7012 13948 7064 14000
rect 7380 13991 7432 14000
rect 7380 13957 7389 13991
rect 7389 13957 7423 13991
rect 7423 13957 7432 13991
rect 7380 13948 7432 13957
rect 9680 13948 9732 14000
rect 9772 13948 9824 14000
rect 3976 13880 4028 13932
rect 9956 13923 10008 13932
rect 2044 13812 2096 13864
rect 4528 13855 4580 13864
rect 4528 13821 4537 13855
rect 4537 13821 4571 13855
rect 4571 13821 4580 13855
rect 4528 13812 4580 13821
rect 4620 13812 4672 13864
rect 6000 13855 6052 13864
rect 6000 13821 6009 13855
rect 6009 13821 6043 13855
rect 6043 13821 6052 13855
rect 6000 13812 6052 13821
rect 6644 13787 6696 13796
rect 6644 13753 6653 13787
rect 6653 13753 6687 13787
rect 6687 13753 6696 13787
rect 6644 13744 6696 13753
rect 6920 13812 6972 13864
rect 3516 13676 3568 13728
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 10416 13880 10468 13932
rect 11980 14016 12032 14068
rect 14372 14016 14424 14068
rect 22468 14016 22520 14068
rect 12808 13991 12860 14000
rect 12808 13957 12817 13991
rect 12817 13957 12851 13991
rect 12851 13957 12860 13991
rect 12808 13948 12860 13957
rect 14280 13991 14332 14000
rect 14280 13957 14289 13991
rect 14289 13957 14323 13991
rect 14323 13957 14332 13991
rect 14280 13948 14332 13957
rect 14832 13991 14884 14000
rect 14832 13957 14841 13991
rect 14841 13957 14875 13991
rect 14875 13957 14884 13991
rect 14832 13948 14884 13957
rect 15476 13991 15528 14000
rect 15476 13957 15485 13991
rect 15485 13957 15519 13991
rect 15519 13957 15528 13991
rect 15476 13948 15528 13957
rect 15568 13948 15620 14000
rect 17684 13880 17736 13932
rect 17868 13880 17920 13932
rect 18420 13880 18472 13932
rect 19984 13948 20036 14000
rect 22100 13991 22152 14000
rect 18788 13880 18840 13932
rect 20996 13923 21048 13932
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 12256 13812 12308 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 15108 13812 15160 13864
rect 17408 13812 17460 13864
rect 20168 13812 20220 13864
rect 22100 13957 22109 13991
rect 22109 13957 22143 13991
rect 22143 13957 22152 13991
rect 22100 13948 22152 13957
rect 23480 13948 23532 14000
rect 32404 13948 32456 14000
rect 22744 13923 22796 13932
rect 22744 13889 22753 13923
rect 22753 13889 22787 13923
rect 22787 13889 22796 13923
rect 23388 13923 23440 13932
rect 22744 13880 22796 13889
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 22468 13812 22520 13864
rect 9404 13744 9456 13796
rect 9496 13744 9548 13796
rect 12900 13744 12952 13796
rect 19248 13744 19300 13796
rect 10600 13676 10652 13728
rect 11152 13676 11204 13728
rect 18972 13676 19024 13728
rect 19156 13719 19208 13728
rect 19156 13685 19165 13719
rect 19165 13685 19199 13719
rect 19199 13685 19208 13719
rect 19156 13676 19208 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1952 13472 2004 13524
rect 2412 13472 2464 13524
rect 4712 13472 4764 13524
rect 4988 13472 5040 13524
rect 4804 13404 4856 13456
rect 5448 13404 5500 13456
rect 6644 13472 6696 13524
rect 8852 13472 8904 13524
rect 9128 13472 9180 13524
rect 9220 13472 9272 13524
rect 14280 13472 14332 13524
rect 15384 13472 15436 13524
rect 15476 13472 15528 13524
rect 17960 13472 18012 13524
rect 18788 13472 18840 13524
rect 20076 13472 20128 13524
rect 21640 13472 21692 13524
rect 22468 13515 22520 13524
rect 22468 13481 22477 13515
rect 22477 13481 22511 13515
rect 22511 13481 22520 13515
rect 22468 13472 22520 13481
rect 6460 13336 6512 13388
rect 8116 13404 8168 13456
rect 13544 13404 13596 13456
rect 15292 13404 15344 13456
rect 18972 13404 19024 13456
rect 20812 13447 20864 13456
rect 20812 13413 20821 13447
rect 20821 13413 20855 13447
rect 20855 13413 20864 13447
rect 20812 13404 20864 13413
rect 20996 13404 21048 13456
rect 5356 13268 5408 13320
rect 5540 13268 5592 13320
rect 5632 13268 5684 13320
rect 8668 13336 8720 13388
rect 11152 13336 11204 13388
rect 6000 13200 6052 13252
rect 9956 13268 10008 13320
rect 10416 13268 10468 13320
rect 11336 13268 11388 13320
rect 11520 13268 11572 13320
rect 13452 13268 13504 13320
rect 13820 13268 13872 13320
rect 16764 13336 16816 13388
rect 20904 13336 20956 13388
rect 18788 13311 18840 13320
rect 18788 13277 18797 13311
rect 18797 13277 18831 13311
rect 18831 13277 18840 13311
rect 18788 13268 18840 13277
rect 19984 13268 20036 13320
rect 22192 13268 22244 13320
rect 23388 13268 23440 13320
rect 35900 13311 35952 13320
rect 35900 13277 35909 13311
rect 35909 13277 35943 13311
rect 35943 13277 35952 13311
rect 35900 13268 35952 13277
rect 6460 13132 6512 13184
rect 6828 13243 6880 13252
rect 6828 13209 6837 13243
rect 6837 13209 6871 13243
rect 6871 13209 6880 13243
rect 6828 13200 6880 13209
rect 7104 13200 7156 13252
rect 9128 13243 9180 13252
rect 9128 13209 9137 13243
rect 9137 13209 9171 13243
rect 9171 13209 9180 13243
rect 9128 13200 9180 13209
rect 12164 13243 12216 13252
rect 12164 13209 12173 13243
rect 12173 13209 12207 13243
rect 12207 13209 12216 13243
rect 12164 13200 12216 13209
rect 9956 13132 10008 13184
rect 13176 13200 13228 13252
rect 13728 13200 13780 13252
rect 12348 13132 12400 13184
rect 14924 13200 14976 13252
rect 17224 13200 17276 13252
rect 17408 13243 17460 13252
rect 17408 13209 17417 13243
rect 17417 13209 17451 13243
rect 17451 13209 17460 13243
rect 17408 13200 17460 13209
rect 36084 13175 36136 13184
rect 36084 13141 36093 13175
rect 36093 13141 36127 13175
rect 36127 13141 36136 13175
rect 36084 13132 36136 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 2964 12928 3016 12980
rect 2872 12860 2924 12912
rect 4620 12860 4672 12912
rect 7748 12928 7800 12980
rect 7932 12928 7984 12980
rect 3976 12792 4028 12844
rect 5448 12792 5500 12844
rect 6736 12792 6788 12844
rect 9496 12928 9548 12980
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 10508 12928 10560 12980
rect 12808 12928 12860 12980
rect 12900 12928 12952 12980
rect 9404 12860 9456 12912
rect 13176 12903 13228 12912
rect 9956 12792 10008 12844
rect 13176 12869 13185 12903
rect 13185 12869 13219 12903
rect 13219 12869 13228 12903
rect 13176 12860 13228 12869
rect 14372 12903 14424 12912
rect 14372 12869 14381 12903
rect 14381 12869 14415 12903
rect 14415 12869 14424 12903
rect 14372 12860 14424 12869
rect 2320 12724 2372 12776
rect 3700 12724 3752 12776
rect 4712 12724 4764 12776
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 8208 12724 8260 12776
rect 9496 12724 9548 12776
rect 5724 12656 5776 12708
rect 8668 12656 8720 12708
rect 14004 12724 14056 12776
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 12992 12656 13044 12708
rect 13360 12656 13412 12708
rect 3608 12588 3660 12640
rect 6552 12588 6604 12640
rect 13728 12656 13780 12708
rect 15384 12588 15436 12640
rect 17408 12928 17460 12980
rect 22192 12928 22244 12980
rect 16672 12860 16724 12912
rect 19156 12860 19208 12912
rect 19432 12903 19484 12912
rect 19432 12869 19441 12903
rect 19441 12869 19475 12903
rect 19475 12869 19484 12903
rect 19432 12860 19484 12869
rect 20260 12860 20312 12912
rect 20536 12860 20588 12912
rect 18328 12792 18380 12844
rect 19984 12792 20036 12844
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 18144 12724 18196 12776
rect 19248 12767 19300 12776
rect 19248 12733 19257 12767
rect 19257 12733 19291 12767
rect 19291 12733 19300 12767
rect 19248 12724 19300 12733
rect 16580 12656 16632 12708
rect 35808 12792 35860 12844
rect 22100 12656 22152 12708
rect 18788 12588 18840 12640
rect 18972 12588 19024 12640
rect 20076 12588 20128 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1860 12384 1912 12436
rect 2504 12384 2556 12436
rect 5356 12384 5408 12436
rect 6000 12384 6052 12436
rect 9312 12427 9364 12436
rect 6736 12316 6788 12368
rect 9312 12393 9321 12427
rect 9321 12393 9355 12427
rect 9355 12393 9364 12427
rect 9312 12384 9364 12393
rect 9864 12384 9916 12436
rect 10968 12384 11020 12436
rect 13636 12427 13688 12436
rect 13636 12393 13645 12427
rect 13645 12393 13679 12427
rect 13679 12393 13688 12427
rect 13636 12384 13688 12393
rect 14372 12427 14424 12436
rect 14372 12393 14381 12427
rect 14381 12393 14415 12427
rect 14415 12393 14424 12427
rect 14372 12384 14424 12393
rect 3976 12180 4028 12232
rect 6920 12248 6972 12300
rect 7288 12248 7340 12300
rect 8668 12248 8720 12300
rect 9864 12248 9916 12300
rect 6368 12180 6420 12232
rect 6828 12180 6880 12232
rect 8760 12180 8812 12232
rect 9496 12180 9548 12232
rect 9772 12180 9824 12232
rect 9956 12180 10008 12232
rect 10692 12180 10744 12232
rect 11612 12248 11664 12300
rect 11704 12248 11756 12300
rect 5356 12044 5408 12096
rect 5724 12155 5776 12164
rect 5724 12121 5733 12155
rect 5733 12121 5767 12155
rect 5767 12121 5776 12155
rect 5724 12112 5776 12121
rect 6920 12044 6972 12096
rect 8024 12044 8076 12096
rect 8392 12112 8444 12164
rect 8668 12112 8720 12164
rect 11428 12112 11480 12164
rect 14004 12316 14056 12368
rect 15936 12384 15988 12436
rect 16672 12427 16724 12436
rect 16672 12393 16681 12427
rect 16681 12393 16715 12427
rect 16715 12393 16724 12427
rect 16672 12384 16724 12393
rect 16856 12384 16908 12436
rect 12072 12248 12124 12300
rect 17408 12316 17460 12368
rect 18972 12384 19024 12436
rect 16580 12248 16632 12300
rect 35532 12248 35584 12300
rect 14464 12223 14516 12232
rect 12992 12155 13044 12164
rect 9312 12044 9364 12096
rect 10968 12044 11020 12096
rect 12992 12121 13001 12155
rect 13001 12121 13035 12155
rect 13035 12121 13044 12155
rect 12992 12112 13044 12121
rect 11796 12044 11848 12096
rect 14004 12044 14056 12096
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 16764 12223 16816 12232
rect 16764 12189 16773 12223
rect 16773 12189 16807 12223
rect 16807 12189 16816 12223
rect 16764 12180 16816 12189
rect 15476 12155 15528 12164
rect 15476 12121 15485 12155
rect 15485 12121 15519 12155
rect 15519 12121 15528 12155
rect 15476 12112 15528 12121
rect 15568 12112 15620 12164
rect 15660 12044 15712 12096
rect 15936 12044 15988 12096
rect 17592 12044 17644 12096
rect 17776 12155 17828 12164
rect 17776 12121 17792 12155
rect 17792 12121 17826 12155
rect 17826 12121 17828 12155
rect 17776 12112 17828 12121
rect 20076 12155 20128 12164
rect 20076 12121 20085 12155
rect 20085 12121 20119 12155
rect 20119 12121 20128 12155
rect 20076 12112 20128 12121
rect 21088 12044 21140 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 1676 11840 1728 11892
rect 1768 11840 1820 11892
rect 3332 11772 3384 11824
rect 7564 11840 7616 11892
rect 10048 11883 10100 11892
rect 3884 11636 3936 11688
rect 3516 11568 3568 11620
rect 1676 11500 1728 11552
rect 4712 11636 4764 11688
rect 4988 11636 5040 11688
rect 5356 11568 5408 11620
rect 7840 11772 7892 11824
rect 8300 11772 8352 11824
rect 10048 11849 10057 11883
rect 10057 11849 10091 11883
rect 10091 11849 10100 11883
rect 10048 11840 10100 11849
rect 10324 11772 10376 11824
rect 10876 11815 10928 11824
rect 10876 11781 10885 11815
rect 10885 11781 10919 11815
rect 10919 11781 10928 11815
rect 10876 11772 10928 11781
rect 11428 11772 11480 11824
rect 13176 11840 13228 11892
rect 15476 11840 15528 11892
rect 16212 11840 16264 11892
rect 6276 11704 6328 11756
rect 6828 11704 6880 11756
rect 10232 11747 10284 11756
rect 10232 11713 10241 11747
rect 10241 11713 10275 11747
rect 10275 11713 10284 11747
rect 10232 11704 10284 11713
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 14004 11704 14056 11756
rect 14464 11704 14516 11756
rect 14556 11704 14608 11756
rect 15200 11704 15252 11756
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 17132 11772 17184 11824
rect 17408 11815 17460 11824
rect 17408 11781 17417 11815
rect 17417 11781 17451 11815
rect 17451 11781 17460 11815
rect 17408 11772 17460 11781
rect 17592 11772 17644 11824
rect 19432 11840 19484 11892
rect 16488 11704 16540 11756
rect 20260 11772 20312 11824
rect 20812 11840 20864 11892
rect 6184 11636 6236 11688
rect 7288 11636 7340 11688
rect 5908 11568 5960 11620
rect 11796 11636 11848 11688
rect 9220 11568 9272 11620
rect 12532 11636 12584 11688
rect 16764 11636 16816 11688
rect 17592 11636 17644 11688
rect 18236 11636 18288 11688
rect 6276 11500 6328 11552
rect 10784 11500 10836 11552
rect 14464 11500 14516 11552
rect 14556 11500 14608 11552
rect 16856 11500 16908 11552
rect 17868 11611 17920 11620
rect 17868 11577 17877 11611
rect 17877 11577 17911 11611
rect 17911 11577 17920 11611
rect 17868 11568 17920 11577
rect 18052 11500 18104 11552
rect 18512 11543 18564 11552
rect 18512 11509 18521 11543
rect 18521 11509 18555 11543
rect 18555 11509 18564 11543
rect 18512 11500 18564 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3608 11296 3660 11348
rect 5172 11296 5224 11348
rect 5724 11296 5776 11348
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 13820 11296 13872 11348
rect 14280 11296 14332 11348
rect 17500 11296 17552 11348
rect 12532 11228 12584 11280
rect 1584 11092 1636 11144
rect 3884 11160 3936 11212
rect 3976 11160 4028 11212
rect 5724 11160 5776 11212
rect 7288 11160 7340 11212
rect 9496 11160 9548 11212
rect 17040 11228 17092 11280
rect 17868 11228 17920 11280
rect 36268 11271 36320 11280
rect 36268 11237 36277 11271
rect 36277 11237 36311 11271
rect 36311 11237 36320 11271
rect 36268 11228 36320 11237
rect 14832 11203 14884 11212
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 11796 11092 11848 11144
rect 12716 11092 12768 11144
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15384 11160 15436 11212
rect 15936 11160 15988 11212
rect 16580 11160 16632 11212
rect 1952 11067 2004 11076
rect 1952 11033 1961 11067
rect 1961 11033 1995 11067
rect 1995 11033 2004 11067
rect 1952 11024 2004 11033
rect 4988 11024 5040 11076
rect 6276 11024 6328 11076
rect 6828 11024 6880 11076
rect 6920 11024 6972 11076
rect 8392 11024 8444 11076
rect 9036 11024 9088 11076
rect 9864 11024 9916 11076
rect 6000 10956 6052 11008
rect 9220 10956 9272 11008
rect 10692 10956 10744 11008
rect 12624 10956 12676 11008
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 14648 11024 14700 11076
rect 15568 10956 15620 11008
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 17500 11024 17552 11076
rect 18052 11067 18104 11076
rect 18052 11033 18061 11067
rect 18061 11033 18095 11067
rect 18095 11033 18104 11067
rect 36084 11135 36136 11144
rect 36084 11101 36093 11135
rect 36093 11101 36127 11135
rect 36127 11101 36136 11135
rect 36084 11092 36136 11101
rect 18052 11024 18104 11033
rect 19340 11024 19392 11076
rect 17592 10956 17644 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3884 10795 3936 10804
rect 3884 10761 3893 10795
rect 3893 10761 3927 10795
rect 3927 10761 3936 10795
rect 3884 10752 3936 10761
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 7472 10752 7524 10804
rect 8484 10684 8536 10736
rect 14556 10752 14608 10804
rect 2688 10616 2740 10668
rect 6828 10659 6880 10668
rect 4804 10548 4856 10600
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 7288 10616 7340 10668
rect 7840 10591 7892 10600
rect 7840 10557 7849 10591
rect 7849 10557 7883 10591
rect 7883 10557 7892 10591
rect 7840 10548 7892 10557
rect 8300 10548 8352 10600
rect 11704 10684 11756 10736
rect 9220 10616 9272 10668
rect 10876 10659 10928 10668
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 14096 10684 14148 10736
rect 14740 10727 14792 10736
rect 14740 10693 14749 10727
rect 14749 10693 14783 10727
rect 14783 10693 14792 10727
rect 14740 10684 14792 10693
rect 17684 10752 17736 10804
rect 15844 10684 15896 10736
rect 18512 10684 18564 10736
rect 13268 10616 13320 10668
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 17592 10659 17644 10668
rect 17592 10625 17601 10659
rect 17601 10625 17635 10659
rect 17635 10625 17644 10659
rect 17592 10616 17644 10625
rect 21824 10752 21876 10804
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 11612 10548 11664 10600
rect 15660 10591 15712 10600
rect 7564 10480 7616 10532
rect 10232 10480 10284 10532
rect 12716 10480 12768 10532
rect 14280 10523 14332 10532
rect 14280 10489 14289 10523
rect 14289 10489 14323 10523
rect 14323 10489 14332 10523
rect 14280 10480 14332 10489
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 16948 10591 17000 10600
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 15752 10480 15804 10532
rect 4896 10455 4948 10464
rect 4896 10421 4905 10455
rect 4905 10421 4939 10455
rect 4939 10421 4948 10455
rect 4896 10412 4948 10421
rect 7288 10412 7340 10464
rect 7932 10412 7984 10464
rect 11980 10412 12032 10464
rect 13176 10412 13228 10464
rect 14832 10412 14884 10464
rect 19432 10412 19484 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 3976 10208 4028 10260
rect 3792 10140 3844 10192
rect 1584 10115 1636 10124
rect 1584 10081 1593 10115
rect 1593 10081 1627 10115
rect 1627 10081 1636 10115
rect 1584 10072 1636 10081
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 4620 10072 4672 10124
rect 4896 10004 4948 10056
rect 8300 10208 8352 10260
rect 8484 10251 8536 10260
rect 8484 10217 8493 10251
rect 8493 10217 8527 10251
rect 8527 10217 8536 10251
rect 8484 10208 8536 10217
rect 11888 10208 11940 10260
rect 15844 10251 15896 10260
rect 7564 10140 7616 10192
rect 10784 10140 10836 10192
rect 15844 10217 15853 10251
rect 15853 10217 15887 10251
rect 15887 10217 15896 10251
rect 15844 10208 15896 10217
rect 5724 10115 5776 10124
rect 5724 10081 5733 10115
rect 5733 10081 5767 10115
rect 5767 10081 5776 10115
rect 5724 10072 5776 10081
rect 6092 10072 6144 10124
rect 9220 10004 9272 10056
rect 10600 10072 10652 10124
rect 11888 10072 11940 10124
rect 12072 10115 12124 10124
rect 12072 10081 12081 10115
rect 12081 10081 12115 10115
rect 12115 10081 12124 10115
rect 12072 10072 12124 10081
rect 13820 10072 13872 10124
rect 18144 10072 18196 10124
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 4804 9868 4856 9920
rect 5264 9868 5316 9920
rect 6092 9936 6144 9988
rect 7012 9936 7064 9988
rect 8484 9936 8536 9988
rect 9772 9936 9824 9988
rect 15200 10004 15252 10056
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 7840 9868 7892 9920
rect 10600 9868 10652 9920
rect 11796 9936 11848 9988
rect 11980 9979 12032 9988
rect 11980 9945 11989 9979
rect 11989 9945 12023 9979
rect 12023 9945 12032 9979
rect 11980 9936 12032 9945
rect 13176 9979 13228 9988
rect 13176 9945 13185 9979
rect 13185 9945 13219 9979
rect 13219 9945 13228 9979
rect 13176 9936 13228 9945
rect 14280 9979 14332 9988
rect 14280 9945 14289 9979
rect 14289 9945 14323 9979
rect 14323 9945 14332 9979
rect 14280 9936 14332 9945
rect 14832 9979 14884 9988
rect 14832 9945 14841 9979
rect 14841 9945 14875 9979
rect 14875 9945 14884 9979
rect 14832 9936 14884 9945
rect 14096 9868 14148 9920
rect 16488 9911 16540 9920
rect 16488 9877 16497 9911
rect 16497 9877 16531 9911
rect 16531 9877 16540 9911
rect 16488 9868 16540 9877
rect 17040 9911 17092 9920
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 17040 9868 17092 9877
rect 35440 9868 35492 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2688 9664 2740 9716
rect 5540 9664 5592 9716
rect 6828 9664 6880 9716
rect 2504 9596 2556 9648
rect 3148 9596 3200 9648
rect 3332 9596 3384 9648
rect 5908 9596 5960 9648
rect 6920 9596 6972 9648
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 8392 9664 8444 9716
rect 9128 9664 9180 9716
rect 8668 9596 8720 9648
rect 8760 9528 8812 9580
rect 9588 9664 9640 9716
rect 9864 9596 9916 9648
rect 12992 9664 13044 9716
rect 16488 9664 16540 9716
rect 17684 9664 17736 9716
rect 36084 9664 36136 9716
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 4896 9460 4948 9512
rect 5172 9460 5224 9512
rect 5264 9460 5316 9512
rect 9404 9460 9456 9512
rect 9680 9460 9732 9512
rect 10048 9460 10100 9512
rect 10324 9528 10376 9580
rect 12072 9596 12124 9648
rect 11980 9528 12032 9580
rect 13084 9528 13136 9580
rect 13820 9528 13872 9580
rect 15016 9596 15068 9648
rect 14556 9528 14608 9580
rect 6552 9392 6604 9444
rect 5540 9324 5592 9376
rect 6092 9324 6144 9376
rect 8852 9392 8904 9444
rect 8300 9324 8352 9376
rect 10508 9392 10560 9444
rect 14648 9460 14700 9512
rect 15108 9528 15160 9580
rect 18604 9460 18656 9512
rect 12992 9392 13044 9444
rect 9864 9324 9916 9376
rect 14280 9392 14332 9444
rect 13176 9324 13228 9376
rect 15476 9324 15528 9376
rect 27160 9324 27212 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 6000 9120 6052 9172
rect 6368 9052 6420 9104
rect 7564 9052 7616 9104
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 8852 9120 8904 9172
rect 9496 9052 9548 9104
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 5264 8984 5316 9036
rect 5724 8984 5776 9036
rect 8392 8984 8444 9036
rect 9864 8984 9916 9036
rect 11060 9120 11112 9172
rect 14832 9120 14884 9172
rect 14924 9163 14976 9172
rect 14924 9129 14933 9163
rect 14933 9129 14967 9163
rect 14967 9129 14976 9163
rect 14924 9120 14976 9129
rect 10048 9052 10100 9104
rect 12440 9052 12492 9104
rect 36084 9095 36136 9104
rect 36084 9061 36093 9095
rect 36093 9061 36127 9095
rect 36127 9061 36136 9095
rect 36084 9052 36136 9061
rect 4620 8916 4672 8968
rect 6552 8916 6604 8968
rect 7472 8916 7524 8968
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 8484 8916 8536 8968
rect 8760 8916 8812 8968
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 10600 8916 10652 8968
rect 14740 8984 14792 9036
rect 1952 8891 2004 8900
rect 1952 8857 1961 8891
rect 1961 8857 1995 8891
rect 1995 8857 2004 8891
rect 1952 8848 2004 8857
rect 2044 8848 2096 8900
rect 6092 8848 6144 8900
rect 6276 8848 6328 8900
rect 6000 8780 6052 8832
rect 7380 8848 7432 8900
rect 12716 8916 12768 8968
rect 16856 8848 16908 8900
rect 36268 8891 36320 8900
rect 36268 8857 36277 8891
rect 36277 8857 36311 8891
rect 36311 8857 36320 8891
rect 36268 8848 36320 8857
rect 12532 8780 12584 8832
rect 15108 8780 15160 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 4896 8576 4948 8628
rect 2688 8508 2740 8560
rect 3424 8508 3476 8560
rect 3608 8508 3660 8560
rect 5540 8508 5592 8560
rect 5816 8576 5868 8628
rect 6460 8576 6512 8628
rect 9312 8619 9364 8628
rect 9312 8585 9321 8619
rect 9321 8585 9355 8619
rect 9355 8585 9364 8619
rect 9312 8576 9364 8585
rect 11336 8576 11388 8628
rect 11704 8576 11756 8628
rect 12440 8576 12492 8628
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 14004 8619 14056 8628
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 14556 8619 14608 8628
rect 14556 8585 14565 8619
rect 14565 8585 14599 8619
rect 14599 8585 14608 8619
rect 14556 8576 14608 8585
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 6276 8508 6328 8560
rect 3884 8440 3936 8492
rect 4896 8440 4948 8492
rect 5356 8440 5408 8492
rect 6736 8440 6788 8492
rect 7288 8440 7340 8492
rect 7472 8440 7524 8492
rect 8484 8483 8536 8492
rect 7748 8372 7800 8424
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 9680 8508 9732 8560
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 10140 8508 10192 8560
rect 10416 8551 10468 8560
rect 10416 8517 10425 8551
rect 10425 8517 10459 8551
rect 10459 8517 10468 8551
rect 10416 8508 10468 8517
rect 11888 8508 11940 8560
rect 9404 8440 9456 8449
rect 9312 8372 9364 8424
rect 11612 8372 11664 8424
rect 2688 8304 2740 8356
rect 18604 8440 18656 8492
rect 3424 8236 3476 8288
rect 7104 8279 7156 8288
rect 7104 8245 7113 8279
rect 7113 8245 7147 8279
rect 7147 8245 7156 8279
rect 7104 8236 7156 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3240 8032 3292 8084
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 6552 8032 6604 8084
rect 7380 8032 7432 8084
rect 10968 8032 11020 8084
rect 5080 7964 5132 8016
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 3056 7828 3108 7880
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 5632 7828 5684 7880
rect 7288 7896 7340 7948
rect 8300 7828 8352 7880
rect 8484 7828 8536 7880
rect 8944 7828 8996 7880
rect 9220 7828 9272 7880
rect 3792 7760 3844 7812
rect 5448 7692 5500 7744
rect 8944 7692 8996 7744
rect 11980 7692 12032 7744
rect 13084 7964 13136 8016
rect 13728 8032 13780 8084
rect 36636 8032 36688 8084
rect 14188 7964 14240 8016
rect 14096 7896 14148 7948
rect 36268 7803 36320 7812
rect 36268 7769 36277 7803
rect 36277 7769 36311 7803
rect 36311 7769 36320 7803
rect 36268 7760 36320 7769
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 3792 7531 3844 7540
rect 3792 7497 3801 7531
rect 3801 7497 3835 7531
rect 3835 7497 3844 7531
rect 3792 7488 3844 7497
rect 2596 7420 2648 7472
rect 2780 7420 2832 7472
rect 3148 7420 3200 7472
rect 3424 7352 3476 7404
rect 5540 7488 5592 7540
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 8116 7488 8168 7540
rect 10416 7488 10468 7540
rect 12256 7488 12308 7540
rect 5264 7420 5316 7472
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 9588 7420 9640 7472
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 5172 7284 5224 7336
rect 5724 7284 5776 7336
rect 1952 7216 2004 7268
rect 3700 7148 3752 7200
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 9772 7352 9824 7404
rect 12992 7352 13044 7404
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 9680 7216 9732 7268
rect 10600 7259 10652 7268
rect 10600 7225 10609 7259
rect 10609 7225 10643 7259
rect 10643 7225 10652 7259
rect 10600 7216 10652 7225
rect 9772 7148 9824 7200
rect 10324 7148 10376 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 8668 6944 8720 6996
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 3424 6808 3476 6860
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 5908 6851 5960 6860
rect 5908 6817 5917 6851
rect 5917 6817 5951 6851
rect 5951 6817 5960 6851
rect 5908 6808 5960 6817
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 10232 6808 10284 6860
rect 10600 6808 10652 6860
rect 3792 6740 3844 6792
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 2964 6672 3016 6724
rect 2596 6604 2648 6656
rect 6184 6740 6236 6792
rect 19340 6740 19392 6792
rect 9404 6672 9456 6724
rect 11888 6672 11940 6724
rect 13176 6715 13228 6724
rect 13176 6681 13185 6715
rect 13185 6681 13219 6715
rect 13219 6681 13228 6715
rect 13176 6672 13228 6681
rect 13268 6715 13320 6724
rect 13268 6681 13277 6715
rect 13277 6681 13311 6715
rect 13311 6681 13320 6715
rect 13268 6672 13320 6681
rect 3608 6604 3660 6656
rect 7656 6604 7708 6656
rect 8208 6604 8260 6656
rect 17224 6604 17276 6656
rect 24676 6604 24728 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 3700 6400 3752 6452
rect 4620 6400 4672 6452
rect 5632 6400 5684 6452
rect 6552 6443 6604 6452
rect 6552 6409 6561 6443
rect 6561 6409 6595 6443
rect 6595 6409 6604 6443
rect 6552 6400 6604 6409
rect 7840 6400 7892 6452
rect 7932 6400 7984 6452
rect 9036 6443 9088 6452
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 9680 6400 9732 6452
rect 13268 6400 13320 6452
rect 17224 6400 17276 6452
rect 36176 6400 36228 6452
rect 3240 6332 3292 6384
rect 7012 6332 7064 6384
rect 7748 6332 7800 6384
rect 2044 6264 2096 6316
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 4068 6264 4120 6316
rect 2596 6196 2648 6248
rect 5356 6264 5408 6316
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 4068 6128 4120 6180
rect 8484 6128 8536 6180
rect 24584 6128 24636 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1768 5856 1820 5908
rect 2872 5856 2924 5908
rect 3148 5856 3200 5908
rect 4804 5856 4856 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 6552 5856 6604 5908
rect 3792 5788 3844 5840
rect 7748 5788 7800 5840
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 9772 5720 9824 5772
rect 3240 5652 3292 5704
rect 4068 5652 4120 5704
rect 2320 5627 2372 5636
rect 2320 5593 2329 5627
rect 2329 5593 2363 5627
rect 2363 5593 2372 5627
rect 2320 5584 2372 5593
rect 3608 5584 3660 5636
rect 12256 5584 12308 5636
rect 35532 5627 35584 5636
rect 35532 5593 35541 5627
rect 35541 5593 35575 5627
rect 35575 5593 35584 5627
rect 35532 5584 35584 5593
rect 36268 5559 36320 5568
rect 36268 5525 36277 5559
rect 36277 5525 36311 5559
rect 36311 5525 36320 5559
rect 36268 5516 36320 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3056 5312 3108 5364
rect 4712 5312 4764 5364
rect 5632 5312 5684 5364
rect 5724 5355 5776 5364
rect 5724 5321 5733 5355
rect 5733 5321 5767 5355
rect 5767 5321 5776 5355
rect 17684 5355 17736 5364
rect 5724 5312 5776 5321
rect 17684 5321 17693 5355
rect 17693 5321 17727 5355
rect 17727 5321 17736 5355
rect 17684 5312 17736 5321
rect 2412 5244 2464 5296
rect 1952 5176 2004 5228
rect 2596 5219 2648 5228
rect 2596 5185 2605 5219
rect 2605 5185 2639 5219
rect 2639 5185 2648 5219
rect 2596 5176 2648 5185
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 6000 5108 6052 5160
rect 6920 5040 6972 5092
rect 1676 5015 1728 5024
rect 1676 4981 1685 5015
rect 1685 4981 1719 5015
rect 1719 4981 1728 5015
rect 1676 4972 1728 4981
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 17500 4972 17552 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2044 4811 2096 4820
rect 2044 4777 2053 4811
rect 2053 4777 2087 4811
rect 2087 4777 2096 4811
rect 2044 4768 2096 4777
rect 2964 4768 3016 4820
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 3516 4768 3568 4820
rect 4896 4768 4948 4820
rect 5632 4768 5684 4820
rect 1952 4607 2004 4616
rect 1952 4573 1961 4607
rect 1961 4573 1995 4607
rect 1995 4573 2004 4607
rect 1952 4564 2004 4573
rect 3240 4564 3292 4616
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 36084 4607 36136 4616
rect 36084 4573 36093 4607
rect 36093 4573 36127 4607
rect 36127 4573 36136 4607
rect 36084 4564 36136 4573
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 36268 4471 36320 4480
rect 36268 4437 36277 4471
rect 36277 4437 36311 4471
rect 36311 4437 36320 4471
rect 36268 4428 36320 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2412 4224 2464 4276
rect 3792 4224 3844 4276
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 2780 4088 2832 4140
rect 3976 4088 4028 4140
rect 25688 4088 25740 4140
rect 4988 4020 5040 4072
rect 36084 3884 36136 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2780 3680 2832 3732
rect 3884 3476 3936 3528
rect 15936 3476 15988 3528
rect 35808 3476 35860 3528
rect 20352 3408 20404 3460
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 20720 3340 20772 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 35440 3179 35492 3188
rect 35440 3145 35449 3179
rect 35449 3145 35483 3179
rect 35483 3145 35492 3179
rect 35440 3136 35492 3145
rect 36176 3179 36228 3188
rect 36176 3145 36185 3179
rect 36185 3145 36219 3179
rect 36219 3145 36228 3179
rect 36176 3136 36228 3145
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 36728 3068 36780 3120
rect 36360 3000 36412 3052
rect 18880 2932 18932 2984
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 7840 2796 7892 2848
rect 20628 2796 20680 2848
rect 27068 2796 27120 2848
rect 30380 2839 30432 2848
rect 30380 2805 30389 2839
rect 30389 2805 30423 2839
rect 30423 2805 30432 2839
rect 30380 2796 30432 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 7288 2592 7340 2644
rect 12992 2635 13044 2644
rect 12992 2601 13001 2635
rect 13001 2601 13035 2635
rect 13035 2601 13044 2635
rect 12992 2592 13044 2601
rect 18604 2592 18656 2644
rect 29828 2635 29880 2644
rect 29828 2601 29837 2635
rect 29837 2601 29871 2635
rect 29871 2601 29880 2635
rect 29828 2592 29880 2601
rect 30564 2635 30616 2644
rect 30564 2601 30573 2635
rect 30573 2601 30607 2635
rect 30607 2601 30616 2635
rect 30564 2592 30616 2601
rect 32404 2635 32456 2644
rect 32404 2601 32413 2635
rect 32413 2601 32447 2635
rect 32447 2601 32456 2635
rect 32404 2592 32456 2601
rect 33784 2592 33836 2644
rect 20 2524 72 2576
rect 11980 2567 12032 2576
rect 11980 2533 11989 2567
rect 11989 2533 12023 2567
rect 12023 2533 12032 2567
rect 11980 2524 12032 2533
rect 19064 2524 19116 2576
rect 7564 2456 7616 2508
rect 23664 2524 23716 2576
rect 27160 2567 27212 2576
rect 27160 2533 27169 2567
rect 27169 2533 27203 2567
rect 27203 2533 27212 2567
rect 27160 2524 27212 2533
rect 34520 2524 34572 2576
rect 2688 2388 2740 2440
rect 1308 2252 1360 2304
rect 3240 2252 3292 2304
rect 20628 2456 20680 2508
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 9220 2320 9272 2372
rect 9680 2320 9732 2372
rect 4528 2252 4580 2304
rect 6460 2252 6512 2304
rect 7748 2252 7800 2304
rect 11060 2295 11112 2304
rect 11060 2261 11069 2295
rect 11069 2261 11103 2295
rect 11103 2261 11112 2295
rect 12900 2388 12952 2440
rect 14188 2388 14240 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 24676 2388 24728 2440
rect 30380 2388 30432 2440
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 11060 2252 11112 2261
rect 15108 2252 15160 2304
rect 25688 2320 25740 2372
rect 27068 2320 27120 2372
rect 17408 2252 17460 2304
rect 19340 2252 19392 2304
rect 20628 2252 20680 2304
rect 22560 2252 22612 2304
rect 23848 2252 23900 2304
rect 25780 2252 25832 2304
rect 29000 2252 29052 2304
rect 32220 2320 32272 2372
rect 33508 2320 33560 2372
rect 35440 2252 35492 2304
rect 36360 2295 36412 2304
rect 36360 2261 36369 2295
rect 36369 2261 36403 2295
rect 36403 2261 36412 2295
rect 36360 2252 36412 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 13542 39200 13598 39800
rect 14830 39200 14886 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 676 36174 704 39200
rect 1674 37496 1730 37505
rect 1674 37431 1730 37440
rect 1688 36854 1716 37431
rect 1964 37126 1992 39200
rect 2870 38856 2926 38865
rect 2870 38791 2926 38800
rect 2320 37256 2372 37262
rect 2320 37198 2372 37204
rect 1952 37120 2004 37126
rect 1952 37062 2004 37068
rect 1676 36848 1728 36854
rect 1676 36790 1728 36796
rect 1860 36644 1912 36650
rect 1860 36586 1912 36592
rect 1872 36281 1900 36586
rect 1858 36272 1914 36281
rect 1858 36207 1914 36216
rect 664 36168 716 36174
rect 664 36110 716 36116
rect 1584 35624 1636 35630
rect 1584 35566 1636 35572
rect 1596 35465 1624 35566
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1596 35290 1624 35391
rect 1584 35284 1636 35290
rect 1584 35226 1636 35232
rect 1584 32360 1636 32366
rect 1584 32302 1636 32308
rect 1596 32065 1624 32302
rect 1582 32056 1638 32065
rect 1582 31991 1584 32000
rect 1636 31991 1638 32000
rect 1584 31962 1636 31968
rect 1674 30696 1730 30705
rect 1674 30631 1730 30640
rect 1688 30598 1716 30631
rect 1676 30592 1728 30598
rect 1676 30534 1728 30540
rect 2332 30326 2360 37198
rect 2884 37126 2912 38791
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 2964 37188 3016 37194
rect 2964 37130 3016 37136
rect 2872 37120 2924 37126
rect 2872 37062 2924 37068
rect 2504 36304 2556 36310
rect 2504 36246 2556 36252
rect 2320 30320 2372 30326
rect 2320 30262 2372 30268
rect 1584 29164 1636 29170
rect 1584 29106 1636 29112
rect 1596 28665 1624 29106
rect 1768 29028 1820 29034
rect 1768 28970 1820 28976
rect 1582 28656 1638 28665
rect 1582 28591 1638 28600
rect 1676 27328 1728 27334
rect 1674 27296 1676 27305
rect 1728 27296 1730 27305
rect 1674 27231 1730 27240
rect 1492 26852 1544 26858
rect 1492 26794 1544 26800
rect 1400 24336 1452 24342
rect 1400 24278 1452 24284
rect 1412 18970 1440 24278
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1412 15434 1440 18906
rect 1504 17202 1532 26794
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1584 24064 1636 24070
rect 1584 24006 1636 24012
rect 1596 23905 1624 24006
rect 1582 23896 1638 23905
rect 1582 23831 1638 23840
rect 1596 22642 1624 23831
rect 1688 23594 1716 26318
rect 1780 24274 1808 28970
rect 1860 27872 1912 27878
rect 1860 27814 1912 27820
rect 1872 27470 1900 27814
rect 2516 27470 2544 36246
rect 2688 35624 2740 35630
rect 2688 35566 2740 35572
rect 1860 27464 1912 27470
rect 1858 27432 1860 27441
rect 2504 27464 2556 27470
rect 1912 27432 1914 27441
rect 2504 27406 2556 27412
rect 1858 27367 1914 27376
rect 2320 27328 2372 27334
rect 2320 27270 2372 27276
rect 1952 26784 2004 26790
rect 1952 26726 2004 26732
rect 1860 26512 1912 26518
rect 1860 26454 1912 26460
rect 1768 24268 1820 24274
rect 1768 24210 1820 24216
rect 1676 23588 1728 23594
rect 1676 23530 1728 23536
rect 1688 22778 1716 23530
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1676 21888 1728 21894
rect 1674 21856 1676 21865
rect 1728 21856 1730 21865
rect 1674 21791 1730 21800
rect 1872 21554 1900 26454
rect 1964 24750 1992 26726
rect 2136 25968 2188 25974
rect 2136 25910 2188 25916
rect 2044 25832 2096 25838
rect 2044 25774 2096 25780
rect 2056 25362 2084 25774
rect 2044 25356 2096 25362
rect 2044 25298 2096 25304
rect 1952 24744 2004 24750
rect 1952 24686 2004 24692
rect 2148 24410 2176 25910
rect 2228 24880 2280 24886
rect 2228 24822 2280 24828
rect 2136 24404 2188 24410
rect 2136 24346 2188 24352
rect 1952 24200 2004 24206
rect 1952 24142 2004 24148
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 20505 1716 21286
rect 1860 20800 1912 20806
rect 1860 20742 1912 20748
rect 1674 20496 1730 20505
rect 1674 20431 1730 20440
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1596 17678 1624 19314
rect 1674 18456 1730 18465
rect 1674 18391 1730 18400
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 17270 1624 17614
rect 1688 17338 1716 18391
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1596 16658 1624 17206
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 15570 1624 16594
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 1596 14482 1624 15506
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1688 11898 1716 16730
rect 1780 15178 1808 19994
rect 1872 16794 1900 20742
rect 1964 19310 1992 24142
rect 2240 23866 2268 24822
rect 2228 23860 2280 23866
rect 2228 23802 2280 23808
rect 2044 23656 2096 23662
rect 2044 23598 2096 23604
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18222 1992 19246
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1872 16658 1900 16730
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1780 15150 1900 15178
rect 1872 14006 1900 15150
rect 2056 14482 2084 23598
rect 2332 22030 2360 27270
rect 2516 25974 2544 27406
rect 2700 27402 2728 35566
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2688 27396 2740 27402
rect 2688 27338 2740 27344
rect 2688 26308 2740 26314
rect 2688 26250 2740 26256
rect 2504 25968 2556 25974
rect 2504 25910 2556 25916
rect 2596 25900 2648 25906
rect 2596 25842 2648 25848
rect 2504 25832 2556 25838
rect 2504 25774 2556 25780
rect 2412 25220 2464 25226
rect 2412 25162 2464 25168
rect 2424 23322 2452 25162
rect 2412 23316 2464 23322
rect 2412 23258 2464 23264
rect 2516 23202 2544 25774
rect 2424 23174 2544 23202
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 2424 17746 2452 23174
rect 2504 23112 2556 23118
rect 2504 23054 2556 23060
rect 2516 22137 2544 23054
rect 2502 22128 2558 22137
rect 2502 22063 2558 22072
rect 2608 20058 2636 25842
rect 2700 25838 2728 26250
rect 2688 25832 2740 25838
rect 2688 25774 2740 25780
rect 2792 24818 2820 32302
rect 2976 26994 3004 37130
rect 3252 36582 3280 37198
rect 3896 37126 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5184 37262 5212 39200
rect 7116 37330 7144 39200
rect 7104 37324 7156 37330
rect 7104 37266 7156 37272
rect 4252 37256 4304 37262
rect 4252 37198 4304 37204
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 4264 36922 4292 37198
rect 8404 37126 8432 39200
rect 9404 37256 9456 37262
rect 9404 37198 9456 37204
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 4252 36916 4304 36922
rect 4252 36858 4304 36864
rect 3240 36576 3292 36582
rect 3240 36518 3292 36524
rect 2964 26988 3016 26994
rect 2964 26930 3016 26936
rect 3252 26042 3280 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 5724 31816 5776 31822
rect 5724 31758 5776 31764
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4620 30252 4672 30258
rect 4620 30194 4672 30200
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3608 26376 3660 26382
rect 3608 26318 3660 26324
rect 3240 26036 3292 26042
rect 3240 25978 3292 25984
rect 3516 25696 3568 25702
rect 3516 25638 3568 25644
rect 3528 25498 3556 25638
rect 3516 25492 3568 25498
rect 3516 25434 3568 25440
rect 3332 25288 3384 25294
rect 3146 25256 3202 25265
rect 3332 25230 3384 25236
rect 3146 25191 3202 25200
rect 3160 25158 3188 25191
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 2780 24812 2832 24818
rect 2780 24754 2832 24760
rect 2792 23497 2820 24754
rect 3344 24410 3372 25230
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3252 23594 3280 23802
rect 3240 23588 3292 23594
rect 3240 23530 3292 23536
rect 3516 23588 3568 23594
rect 3516 23530 3568 23536
rect 2778 23488 2834 23497
rect 2778 23423 2834 23432
rect 2792 23118 2820 23423
rect 3528 23322 3556 23530
rect 3516 23316 3568 23322
rect 3516 23258 3568 23264
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2780 22704 2832 22710
rect 2780 22646 2832 22652
rect 2792 22030 2820 22646
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2792 21486 2820 21966
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2792 21146 2820 21422
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2884 21146 2912 21286
rect 2780 21140 2832 21146
rect 2780 21082 2832 21088
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2792 20942 2820 21082
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2792 20602 2820 20878
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2792 19922 2820 20538
rect 2976 20398 3004 23122
rect 3240 22092 3292 22098
rect 3528 22094 3556 23258
rect 3240 22034 3292 22040
rect 3436 22066 3556 22094
rect 3252 21894 3280 22034
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2686 19816 2742 19825
rect 2686 19751 2688 19760
rect 2740 19751 2742 19760
rect 2688 19722 2740 19728
rect 3068 19553 3096 21830
rect 3054 19544 3110 19553
rect 3054 19479 3110 19488
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 2516 18426 2544 19110
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2410 17096 2466 17105
rect 2410 17031 2412 17040
rect 2464 17031 2466 17040
rect 2964 17060 3016 17066
rect 2412 17002 2464 17008
rect 2964 17002 3016 17008
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1860 14000 1912 14006
rect 1860 13942 1912 13948
rect 2056 13870 2084 14418
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10130 1624 11086
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 1596 9518 1624 9551
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1688 9042 1716 11494
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 7954 1716 8978
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1688 6866 1716 7890
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1780 5914 1808 11834
rect 1872 10130 1900 12378
rect 1964 11082 1992 13466
rect 2332 12782 2360 15846
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2424 13530 2452 14418
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2516 12442 2544 15846
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 2608 9674 2636 14758
rect 2700 11801 2728 16050
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2792 13705 2820 15914
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2884 13297 2912 15030
rect 2976 14550 3004 17002
rect 3068 15162 3096 19479
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 2870 13288 2926 13297
rect 2870 13223 2926 13232
rect 2792 12986 3004 13002
rect 2792 12980 3016 12986
rect 2792 12974 2964 12980
rect 2686 11792 2742 11801
rect 2686 11727 2742 11736
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2700 9722 2728 10610
rect 2516 9654 2636 9674
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2504 9648 2636 9654
rect 2556 9646 2636 9648
rect 2504 9590 2556 9596
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 1964 8809 1992 8842
rect 1950 8800 2006 8809
rect 1950 8735 2006 8744
rect 1964 7274 1992 8735
rect 2056 8634 2084 8842
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2700 8566 2728 9658
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 2608 6662 2636 7414
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4865 1716 4966
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 1964 4622 1992 5170
rect 2056 4826 2084 6258
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2412 5704 2464 5710
rect 2318 5672 2374 5681
rect 2412 5646 2464 5652
rect 2318 5607 2320 5616
rect 2372 5607 2374 5616
rect 2320 5578 2372 5584
rect 2424 5302 2452 5646
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 4146 1992 4558
rect 2424 4282 2452 5238
rect 2608 5234 2636 6190
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1688 3398 1716 3431
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 1688 1465 1716 2790
rect 2700 2446 2728 8298
rect 2792 7478 2820 12974
rect 2964 12922 3016 12928
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2884 12434 2912 12854
rect 2884 12406 3004 12434
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2778 6896 2834 6905
rect 2976 6882 3004 12406
rect 3160 9654 3188 16594
rect 3252 16182 3280 21830
rect 3436 20874 3464 22066
rect 3620 21486 3648 26318
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25430 4660 30194
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 5000 25838 5028 26794
rect 5264 26444 5316 26450
rect 5264 26386 5316 26392
rect 5276 25974 5304 26386
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 4988 25832 5040 25838
rect 4988 25774 5040 25780
rect 4620 25424 4672 25430
rect 4620 25366 4672 25372
rect 3792 25220 3844 25226
rect 3792 25162 3844 25168
rect 3804 24886 3832 25162
rect 4436 25152 4488 25158
rect 4436 25094 4488 25100
rect 3792 24880 3844 24886
rect 3792 24822 3844 24828
rect 3884 24880 3936 24886
rect 3884 24822 3936 24828
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3804 21729 3832 23666
rect 3896 23526 3924 24822
rect 4448 24614 4476 25094
rect 4632 24834 4660 25366
rect 5000 25158 5028 25774
rect 5736 25770 5764 31758
rect 9416 31482 9444 37198
rect 10336 37126 10364 39200
rect 10692 37256 10744 37262
rect 10692 37198 10744 37204
rect 10784 37256 10836 37262
rect 10784 37198 10836 37204
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 10704 36922 10732 37198
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10796 32026 10824 37198
rect 11624 37126 11652 39200
rect 13556 37126 13584 39200
rect 14844 37466 14872 39200
rect 14832 37460 14884 37466
rect 14832 37402 14884 37408
rect 14844 37262 14872 37402
rect 16120 37324 16172 37330
rect 16120 37266 16172 37272
rect 14004 37256 14056 37262
rect 14004 37198 14056 37204
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 11612 37120 11664 37126
rect 11612 37062 11664 37068
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 12256 36848 12308 36854
rect 12256 36790 12308 36796
rect 10876 36780 10928 36786
rect 10876 36722 10928 36728
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10888 31822 10916 36722
rect 10692 31816 10744 31822
rect 10692 31758 10744 31764
rect 10876 31816 10928 31822
rect 10876 31758 10928 31764
rect 9404 31476 9456 31482
rect 9404 31418 9456 31424
rect 5908 27124 5960 27130
rect 5908 27066 5960 27072
rect 5724 25764 5776 25770
rect 5724 25706 5776 25712
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 4988 25152 5040 25158
rect 4988 25094 5040 25100
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 4540 24806 4660 24834
rect 4540 24682 4568 24806
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 4528 24676 4580 24682
rect 4528 24618 4580 24624
rect 4436 24608 4488 24614
rect 4436 24550 4488 24556
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3884 22976 3936 22982
rect 3884 22918 3936 22924
rect 3896 22094 3924 22918
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3896 22066 4016 22094
rect 3790 21720 3846 21729
rect 3790 21655 3846 21664
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3424 20868 3476 20874
rect 3424 20810 3476 20816
rect 3422 20632 3478 20641
rect 3422 20567 3424 20576
rect 3476 20567 3478 20576
rect 3424 20538 3476 20544
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3344 16794 3372 20334
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3528 19446 3556 19994
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3436 18222 3464 18362
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3514 18184 3570 18193
rect 3514 18119 3570 18128
rect 3528 17814 3556 18119
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3330 13016 3386 13025
rect 3330 12951 3386 12960
rect 3344 11830 3372 12951
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2778 6831 2834 6840
rect 2884 6854 3004 6882
rect 2792 4146 2820 6831
rect 2884 5914 2912 6854
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2976 4826 3004 6666
rect 3068 5370 3096 7822
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3160 5914 3188 7414
rect 3252 6390 3280 8026
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3252 5234 3280 5646
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3252 4622 3280 5170
rect 3344 4826 3372 9590
rect 3436 8566 3464 15030
rect 3528 14278 3556 17750
rect 3620 14618 3648 21422
rect 3882 20632 3938 20641
rect 3882 20567 3938 20576
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3712 14498 3740 17070
rect 3804 15094 3832 17206
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3896 14890 3924 20567
rect 3988 17338 4016 22066
rect 4632 21536 4660 24006
rect 4816 23594 4844 24550
rect 4908 24274 4936 24550
rect 4896 24268 4948 24274
rect 4896 24210 4948 24216
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4896 23044 4948 23050
rect 4896 22986 4948 22992
rect 4908 22642 4936 22986
rect 5000 22778 5028 24686
rect 5080 24200 5132 24206
rect 5080 24142 5132 24148
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4896 22500 4948 22506
rect 4896 22442 4948 22448
rect 4632 21508 4752 21536
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4252 20868 4304 20874
rect 4252 20810 4304 20816
rect 4264 20534 4292 20810
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4080 19378 4108 19858
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4080 18834 4108 19314
rect 4528 19304 4580 19310
rect 4526 19272 4528 19281
rect 4580 19272 4582 19281
rect 4526 19207 4582 19216
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4344 18352 4396 18358
rect 4632 18340 4660 21354
rect 4724 20233 4752 21508
rect 4710 20224 4766 20233
rect 4710 20159 4766 20168
rect 4396 18312 4660 18340
rect 4344 18294 4396 18300
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3988 16658 4016 17070
rect 4080 16794 4108 17682
rect 4448 16998 4476 17682
rect 4724 17610 4752 20159
rect 4908 19922 4936 22442
rect 5000 22234 5028 22714
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 5092 21978 5120 24142
rect 5000 21950 5120 21978
rect 5000 21894 5028 21950
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 21010 5028 21830
rect 4988 21004 5040 21010
rect 4988 20946 5040 20952
rect 5080 21004 5132 21010
rect 5080 20946 5132 20952
rect 5092 20890 5120 20946
rect 5184 20913 5212 25094
rect 5264 24268 5316 24274
rect 5264 24210 5316 24216
rect 5276 22506 5304 24210
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 5368 23662 5396 24006
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5460 23526 5488 25094
rect 5552 24886 5580 25230
rect 5540 24880 5592 24886
rect 5540 24822 5592 24828
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5264 22500 5316 22506
rect 5264 22442 5316 22448
rect 5264 21956 5316 21962
rect 5264 21898 5316 21904
rect 5000 20862 5120 20890
rect 5170 20904 5226 20913
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4908 19174 4936 19858
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 5000 18612 5028 20862
rect 5170 20839 5226 20848
rect 5184 19768 5212 20839
rect 5092 19740 5212 19768
rect 5092 18714 5120 19740
rect 5276 19310 5304 21898
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5170 18864 5226 18873
rect 5170 18799 5172 18808
rect 5224 18799 5226 18808
rect 5172 18770 5224 18776
rect 5092 18686 5212 18714
rect 5276 18698 5304 19110
rect 5000 18584 5120 18612
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4250 16688 4306 16697
rect 3976 16652 4028 16658
rect 4724 16658 4752 16934
rect 4250 16623 4252 16632
rect 3976 16594 4028 16600
rect 4304 16623 4306 16632
rect 4712 16652 4764 16658
rect 4252 16594 4304 16600
rect 4712 16594 4764 16600
rect 4724 16561 4752 16594
rect 4710 16552 4766 16561
rect 4710 16487 4766 16496
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4540 16046 4568 16390
rect 4710 16280 4766 16289
rect 4710 16215 4766 16224
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4066 15056 4122 15065
rect 4066 14991 4068 15000
rect 4120 14991 4122 15000
rect 4068 14962 4120 14968
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3620 14470 3740 14498
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3528 11626 3556 13670
rect 3620 12646 3648 14470
rect 3988 14074 4016 14894
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3988 13938 4016 14010
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3988 12850 4016 13874
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3700 12776 3752 12782
rect 3988 12730 4016 12786
rect 3700 12718 3752 12724
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 8090 3464 8230
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3436 6866 3464 7346
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6322 3464 6802
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3528 4826 3556 11562
rect 3620 11354 3648 12582
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3620 6662 3648 8502
rect 3712 7206 3740 12718
rect 3896 12702 4016 12730
rect 3896 11694 3924 12702
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3884 11688 3936 11694
rect 3790 11656 3846 11665
rect 3884 11630 3936 11636
rect 3790 11591 3846 11600
rect 3804 10198 3832 11591
rect 3896 11218 3924 11630
rect 3988 11218 4016 12174
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3896 10810 3924 11154
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3974 10296 4030 10305
rect 3974 10231 3976 10240
rect 4028 10231 4030 10240
rect 3976 10202 4028 10208
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 3804 7546 3832 7754
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 5642 3648 6598
rect 3712 6458 3740 7142
rect 3792 6792 3844 6798
rect 3896 6780 3924 8434
rect 3974 8256 4030 8265
rect 3974 8191 4030 8200
rect 3988 7886 4016 8191
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3844 6752 3924 6780
rect 3792 6734 3844 6740
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3804 5846 3832 6734
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3804 4282 3832 5782
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2792 3738 2820 4082
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3896 3534 3924 4966
rect 3988 4146 4016 7822
rect 4080 6866 4108 14962
rect 4172 14958 4200 15438
rect 4724 15366 4752 16215
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 13870 4568 14214
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 12918 4660 13806
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10130 4660 12854
rect 4724 12782 4752 13466
rect 4816 13462 4844 17478
rect 4986 16552 5042 16561
rect 4896 16516 4948 16522
rect 5092 16522 5120 18584
rect 4986 16487 5042 16496
rect 5080 16516 5132 16522
rect 4896 16458 4948 16464
rect 4908 16250 4936 16458
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 5000 16114 5028 16487
rect 5080 16458 5132 16464
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4908 12594 4936 15302
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4724 12566 4936 12594
rect 4724 12434 4752 12566
rect 4724 12406 4844 12434
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4632 6458 4660 8910
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4080 6186 4108 6258
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5710 4108 6122
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4724 5370 4752 11630
rect 4816 10606 4844 12406
rect 5000 11694 5028 13466
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10062 4936 10406
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 5914 4844 9862
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 8634 4936 9454
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4894 8528 4950 8537
rect 4894 8463 4896 8472
rect 4948 8463 4950 8472
rect 4896 8434 4948 8440
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4908 4826 4936 8434
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 5000 4078 5028 11018
rect 5092 8022 5120 16458
rect 5184 16454 5212 18686
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5262 18320 5318 18329
rect 5262 18255 5318 18264
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5276 16289 5304 18255
rect 5368 16454 5396 20470
rect 5460 18329 5488 21422
rect 5552 20534 5580 22918
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5552 19514 5580 20470
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5552 18426 5580 19178
rect 5644 19009 5672 24754
rect 5736 23662 5764 25706
rect 5816 25220 5868 25226
rect 5816 25162 5868 25168
rect 5828 24410 5856 25162
rect 5920 24818 5948 27066
rect 8576 27056 8628 27062
rect 8576 26998 8628 27004
rect 7932 26920 7984 26926
rect 7932 26862 7984 26868
rect 6736 26580 6788 26586
rect 6736 26522 6788 26528
rect 6644 24880 6696 24886
rect 6644 24822 6696 24828
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 6184 24676 6236 24682
rect 6184 24618 6236 24624
rect 6368 24676 6420 24682
rect 6368 24618 6420 24624
rect 5816 24404 5868 24410
rect 5816 24346 5868 24352
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 5828 23474 5856 23802
rect 5736 23446 5856 23474
rect 5736 19530 5764 23446
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 5828 20992 5856 23258
rect 6000 22704 6052 22710
rect 6000 22646 6052 22652
rect 6012 21060 6040 22646
rect 6196 21978 6224 24618
rect 6380 23322 6408 24618
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6368 23316 6420 23322
rect 6368 23258 6420 23264
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6288 22710 6316 22918
rect 6276 22704 6328 22710
rect 6276 22646 6328 22652
rect 6472 22094 6500 23802
rect 6552 22500 6604 22506
rect 6552 22442 6604 22448
rect 6380 22066 6500 22094
rect 6196 21950 6316 21978
rect 6012 21032 6224 21060
rect 5828 20964 6132 20992
rect 6000 20868 6052 20874
rect 6000 20810 6052 20816
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5920 19922 5948 20334
rect 5908 19916 5960 19922
rect 5908 19858 5960 19864
rect 5736 19514 5856 19530
rect 5736 19508 5868 19514
rect 5736 19502 5816 19508
rect 5736 19334 5764 19502
rect 5816 19450 5868 19456
rect 5736 19306 5856 19334
rect 5630 19000 5686 19009
rect 5828 18986 5856 19306
rect 5630 18935 5686 18944
rect 5736 18958 5856 18986
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5446 18320 5502 18329
rect 5644 18306 5672 18770
rect 5446 18255 5502 18264
rect 5552 18278 5672 18306
rect 5552 17338 5580 18278
rect 5632 18216 5684 18222
rect 5736 18204 5764 18958
rect 5920 18290 5948 19858
rect 6012 18426 6040 20810
rect 6104 18970 6132 20964
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5684 18176 5764 18204
rect 5632 18158 5684 18164
rect 6196 18086 6224 21032
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 5724 17536 5776 17542
rect 5776 17484 5948 17490
rect 5724 17478 5948 17484
rect 5736 17462 5948 17478
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5262 16280 5318 16289
rect 5262 16215 5318 16224
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5184 14074 5212 15982
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5276 14346 5304 15914
rect 5368 15162 5396 16390
rect 5552 16114 5580 16934
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5736 16114 5764 16458
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5368 14414 5396 15098
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5368 13326 5396 14350
rect 5448 13456 5500 13462
rect 5500 13404 5672 13410
rect 5448 13398 5672 13404
rect 5460 13382 5672 13398
rect 5644 13326 5672 13382
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5368 12345 5396 12378
rect 5354 12336 5410 12345
rect 5276 12294 5354 12322
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5184 9518 5212 11290
rect 5276 9926 5304 12294
rect 5354 12271 5410 12280
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11626 5396 12038
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5276 9042 5304 9454
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5368 8616 5396 11562
rect 5184 8588 5396 8616
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5184 7342 5212 8588
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5276 6866 5304 7414
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5368 6798 5396 8434
rect 5460 7750 5488 12786
rect 5552 9722 5580 13262
rect 5736 12714 5764 14486
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11354 5764 12106
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5736 10130 5764 11154
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5552 9466 5580 9658
rect 5552 9438 5672 9466
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 8566 5580 9318
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5552 7546 5580 8502
rect 5644 7886 5672 9438
rect 5736 9042 5764 10066
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5736 8090 5764 8978
rect 5828 8634 5856 14214
rect 5920 11626 5948 17462
rect 6288 17320 6316 21950
rect 6380 18902 6408 22066
rect 6564 21962 6592 22442
rect 6552 21956 6604 21962
rect 6552 21898 6604 21904
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6472 21010 6500 21830
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6472 20534 6500 20810
rect 6460 20528 6512 20534
rect 6460 20470 6512 20476
rect 6564 20398 6592 20878
rect 6656 20777 6684 24822
rect 6748 24750 6776 26522
rect 7944 26450 7972 26862
rect 8208 26512 8260 26518
rect 8208 26454 8260 26460
rect 7932 26444 7984 26450
rect 7932 26386 7984 26392
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 6736 24744 6788 24750
rect 6736 24686 6788 24692
rect 6736 24200 6788 24206
rect 6736 24142 6788 24148
rect 6642 20768 6698 20777
rect 6642 20703 6698 20712
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6472 19514 6500 19654
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6656 18714 6684 20703
rect 6748 20262 6776 24142
rect 6840 23798 6868 25638
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 7024 24410 7052 25162
rect 7944 24886 7972 25638
rect 8220 25430 8248 26454
rect 8588 26042 8616 26998
rect 9220 26852 9272 26858
rect 9220 26794 9272 26800
rect 10600 26852 10652 26858
rect 10600 26794 10652 26800
rect 9232 26450 9260 26794
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 9220 26444 9272 26450
rect 9220 26386 9272 26392
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9784 26042 9812 26250
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 8312 25430 8340 25978
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 8208 25424 8260 25430
rect 8208 25366 8260 25372
rect 8300 25424 8352 25430
rect 8300 25366 8352 25372
rect 8208 25220 8260 25226
rect 8208 25162 8260 25168
rect 7288 24880 7340 24886
rect 7288 24822 7340 24828
rect 7932 24880 7984 24886
rect 7932 24822 7984 24828
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 7116 24206 7144 24346
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7116 23866 7144 24142
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 6828 23792 6880 23798
rect 6828 23734 6880 23740
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 6826 21856 6882 21865
rect 6826 21791 6882 21800
rect 6840 21690 6868 21791
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6840 21010 6868 21422
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 6840 20534 6868 20946
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6748 19786 6776 20198
rect 6828 20052 6880 20058
rect 6932 20040 6960 20470
rect 6880 20012 6960 20040
rect 6828 19994 6880 20000
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 6826 19680 6882 19689
rect 6826 19615 6882 19624
rect 6734 19000 6790 19009
rect 6734 18935 6790 18944
rect 6380 18686 6684 18714
rect 6380 17746 6408 18686
rect 6748 17814 6776 18935
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6196 17292 6316 17320
rect 6000 17196 6052 17202
rect 6196 17184 6224 17292
rect 6052 17156 6224 17184
rect 6276 17196 6328 17202
rect 6000 17138 6052 17144
rect 6276 17138 6328 17144
rect 6012 17105 6040 17138
rect 5998 17096 6054 17105
rect 5998 17031 6054 17040
rect 6012 16697 6040 17031
rect 5998 16688 6054 16697
rect 5998 16623 6054 16632
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 6012 13258 6040 13806
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 6012 12442 6040 13194
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5908 11620 5960 11626
rect 5908 11562 5960 11568
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5552 7410 5580 7482
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 6322 5396 6734
rect 5644 6458 5672 7822
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5644 5370 5672 6394
rect 5736 5370 5764 7278
rect 5920 6866 5948 9590
rect 6012 9178 6040 10950
rect 6104 10130 6132 15370
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 6196 11694 6224 14486
rect 6288 11762 6316 17138
rect 6380 15502 6408 17682
rect 6472 15706 6500 17682
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6656 17338 6684 17546
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6840 17202 6868 19615
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6748 16182 6776 16526
rect 6932 16250 6960 19314
rect 7024 19242 7052 23666
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7208 22574 7236 22986
rect 7300 22710 7328 24822
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 8116 24812 8168 24818
rect 8116 24754 8168 24760
rect 7288 22704 7340 22710
rect 7288 22646 7340 22652
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 7196 22568 7248 22574
rect 7196 22510 7248 22516
rect 7116 22234 7144 22510
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 7116 19378 7144 22170
rect 7208 22098 7236 22510
rect 7392 22438 7420 24754
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 7840 24200 7892 24206
rect 7838 24168 7840 24177
rect 7892 24168 7894 24177
rect 7838 24103 7894 24112
rect 8036 23662 8064 24550
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 8128 23338 8156 24754
rect 8220 24698 8248 25162
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8220 24670 8524 24698
rect 8680 24682 8708 24754
rect 8496 24070 8524 24670
rect 8668 24676 8720 24682
rect 8668 24618 8720 24624
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 7852 23310 8156 23338
rect 7746 23216 7802 23225
rect 7746 23151 7748 23160
rect 7800 23151 7802 23160
rect 7748 23122 7800 23128
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 7196 22092 7248 22098
rect 7196 22034 7248 22040
rect 7208 21486 7236 22034
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7208 20398 7236 21422
rect 7484 20534 7512 22578
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7562 21720 7618 21729
rect 7562 21655 7618 21664
rect 7576 21622 7604 21655
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7196 20392 7248 20398
rect 7576 20380 7604 21558
rect 7668 21185 7696 21966
rect 7654 21176 7710 21185
rect 7654 21111 7710 21120
rect 7196 20334 7248 20340
rect 7392 20352 7604 20380
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 7104 19236 7156 19242
rect 7104 19178 7156 19184
rect 7024 18970 7052 19178
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7116 18873 7144 19178
rect 7208 18970 7236 19246
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7102 18864 7158 18873
rect 7300 18834 7328 19246
rect 7392 19242 7420 20352
rect 7470 20088 7526 20097
rect 7470 20023 7526 20032
rect 7564 20052 7616 20058
rect 7484 19446 7512 20023
rect 7564 19994 7616 20000
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7102 18799 7158 18808
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 7024 16590 7052 18226
rect 7196 18216 7248 18222
rect 7300 18204 7328 18770
rect 7576 18358 7604 19994
rect 7668 19514 7696 19994
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7564 18352 7616 18358
rect 7564 18294 7616 18300
rect 7248 18176 7328 18204
rect 7196 18158 7248 18164
rect 7208 17592 7236 18158
rect 7760 17746 7788 19858
rect 7852 18698 7880 23310
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 7932 22432 7984 22438
rect 8036 22409 8064 22646
rect 7932 22374 7984 22380
rect 8022 22400 8078 22409
rect 7944 22234 7972 22374
rect 8022 22335 8078 22344
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 8036 19961 8064 22335
rect 8128 22030 8156 22918
rect 8404 22681 8432 23054
rect 8390 22672 8446 22681
rect 8390 22607 8446 22616
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8114 21176 8170 21185
rect 8114 21111 8170 21120
rect 8022 19952 8078 19961
rect 8022 19887 8078 19896
rect 8022 19408 8078 19417
rect 8022 19343 8078 19352
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7288 17604 7340 17610
rect 7208 17564 7288 17592
rect 7288 17546 7340 17552
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 7024 16114 7052 16526
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 6734 15872 6790 15881
rect 6734 15807 6790 15816
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6656 13530 6684 13738
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6458 13424 6514 13433
rect 6458 13359 6460 13368
rect 6512 13359 6514 13368
rect 6460 13330 6512 13336
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6642 13152 6698 13161
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 6104 9382 6132 9930
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6090 8936 6146 8945
rect 6090 8871 6092 8880
rect 6144 8871 6146 8880
rect 6092 8842 6144 8848
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5644 4826 5672 5306
rect 6012 5166 6040 8774
rect 6104 5914 6132 8842
rect 6196 6798 6224 11630
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11082 6316 11494
rect 6380 11257 6408 12174
rect 6366 11248 6422 11257
rect 6366 11183 6422 11192
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6380 9110 6408 11183
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6288 8566 6316 8842
rect 6472 8634 6500 13126
rect 6642 13087 6698 13096
rect 6552 12640 6604 12646
rect 6550 12608 6552 12617
rect 6604 12608 6606 12617
rect 6550 12543 6606 12552
rect 6550 12336 6606 12345
rect 6550 12271 6606 12280
rect 6564 11150 6592 12271
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6564 9450 6592 9522
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6564 8090 6592 8910
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6564 7410 6592 8026
rect 6656 7546 6684 13087
rect 6748 12850 6776 15807
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 14482 6960 14894
rect 7024 14618 7052 15914
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6840 14074 6868 14418
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6932 13870 6960 14418
rect 7116 14362 7144 17206
rect 7300 17134 7328 17546
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7300 15978 7328 17070
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16726 7420 16934
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 16182 7420 16390
rect 7668 16182 7696 17478
rect 7838 17368 7894 17377
rect 7838 17303 7894 17312
rect 7852 17270 7880 17303
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 7656 16176 7708 16182
rect 7656 16118 7708 16124
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7024 14346 7144 14362
rect 7012 14340 7144 14346
rect 7064 14334 7144 14340
rect 7012 14282 7064 14288
rect 7392 14006 7420 15302
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7380 14000 7432 14006
rect 7432 13960 7696 13988
rect 7380 13942 7432 13948
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 13433 6960 13806
rect 6918 13424 6974 13433
rect 6918 13359 6974 13368
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6748 12753 6776 12786
rect 6734 12744 6790 12753
rect 6734 12679 6790 12688
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6748 8498 6776 12310
rect 6840 12238 6868 13194
rect 6932 12306 6960 13359
rect 7024 12434 7052 13942
rect 7470 13288 7526 13297
rect 7104 13252 7156 13258
rect 7470 13223 7526 13232
rect 7104 13194 7156 13200
rect 7116 13161 7144 13194
rect 7102 13152 7158 13161
rect 7102 13087 7158 13096
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7024 12406 7236 12434
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6840 11082 6868 11698
rect 6932 11234 6960 12038
rect 6932 11206 7144 11234
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6932 10810 6960 11018
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6840 9722 6868 10610
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6564 5914 6592 6394
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6932 5098 6960 9590
rect 7024 6390 7052 9930
rect 7116 8537 7144 11206
rect 7208 9353 7236 12406
rect 7300 12306 7328 12718
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7300 11694 7328 12242
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7300 11218 7328 11630
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7300 10674 7328 11154
rect 7484 10810 7512 13223
rect 7562 11928 7618 11937
rect 7562 11863 7564 11872
rect 7616 11863 7618 11872
rect 7564 11834 7616 11840
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 9761 7328 10406
rect 7576 10198 7604 10474
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7286 9752 7342 9761
rect 7286 9687 7342 9696
rect 7194 9344 7250 9353
rect 7194 9279 7250 9288
rect 7102 8528 7158 8537
rect 7300 8498 7328 9687
rect 7484 9217 7512 9862
rect 7470 9208 7526 9217
rect 7470 9143 7526 9152
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7392 8809 7420 8842
rect 7378 8800 7434 8809
rect 7378 8735 7434 8744
rect 7484 8673 7512 8910
rect 7470 8664 7526 8673
rect 7470 8599 7526 8608
rect 7102 8463 7158 8472
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7104 8288 7156 8294
rect 7102 8256 7104 8265
rect 7156 8256 7158 8265
rect 7484 8242 7512 8434
rect 7102 8191 7158 8200
rect 7392 8214 7512 8242
rect 7392 8090 7420 8214
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 7300 3058 7328 7890
rect 7470 6896 7526 6905
rect 7470 6831 7472 6840
rect 7524 6831 7526 6840
rect 7472 6802 7524 6808
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7300 2650 7328 2994
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7576 2514 7604 9046
rect 7668 8401 7696 13960
rect 7760 12986 7788 16662
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7760 12050 7788 12922
rect 7852 12434 7880 14282
rect 7944 12986 7972 16526
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7852 12406 7972 12434
rect 7760 12022 7880 12050
rect 7852 11830 7880 12022
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7852 10282 7880 10542
rect 7944 10470 7972 12406
rect 8036 12102 8064 19343
rect 8128 17814 8156 21111
rect 8208 20868 8260 20874
rect 8208 20810 8260 20816
rect 8116 17808 8168 17814
rect 8116 17750 8168 17756
rect 8220 16590 8248 20810
rect 8312 19718 8340 22374
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8404 18714 8432 21082
rect 8496 20058 8524 24006
rect 8668 23588 8720 23594
rect 8668 23530 8720 23536
rect 8574 21992 8630 22001
rect 8574 21927 8630 21936
rect 8588 21894 8616 21927
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8680 21418 8708 23530
rect 8772 21486 8800 25842
rect 8852 25152 8904 25158
rect 8852 25094 8904 25100
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8760 21072 8812 21078
rect 8760 21014 8812 21020
rect 8666 20904 8722 20913
rect 8666 20839 8668 20848
rect 8720 20839 8722 20848
rect 8668 20810 8720 20816
rect 8772 20398 8800 21014
rect 8864 20398 8892 25094
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8956 23798 8984 24550
rect 9232 24342 9260 25842
rect 9692 25294 9720 25910
rect 10520 25838 10548 26726
rect 10612 26518 10640 26794
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10704 26450 10732 31758
rect 12268 30122 12296 36790
rect 14016 36582 14044 37198
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 14004 36576 14056 36582
rect 14004 36518 14056 36524
rect 13820 32836 13872 32842
rect 13820 32778 13872 32784
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 12532 30252 12584 30258
rect 12532 30194 12584 30200
rect 12624 30252 12676 30258
rect 12624 30194 12676 30200
rect 12256 30116 12308 30122
rect 12256 30058 12308 30064
rect 12544 29510 12572 30194
rect 12532 29504 12584 29510
rect 12530 29472 12532 29481
rect 12584 29472 12586 29481
rect 12530 29407 12586 29416
rect 12072 27872 12124 27878
rect 12072 27814 12124 27820
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 11796 27328 11848 27334
rect 11796 27270 11848 27276
rect 11164 26994 11192 27270
rect 11808 27062 11836 27270
rect 11796 27056 11848 27062
rect 11796 26998 11848 27004
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 11152 26988 11204 26994
rect 11152 26930 11204 26936
rect 10968 26784 11020 26790
rect 10968 26726 11020 26732
rect 10692 26444 10744 26450
rect 10692 26386 10744 26392
rect 10980 26314 11008 26726
rect 11900 26586 11928 26998
rect 12084 26926 12112 27814
rect 12636 27606 12664 30194
rect 12624 27600 12676 27606
rect 12624 27542 12676 27548
rect 12072 26920 12124 26926
rect 12072 26862 12124 26868
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 10968 26308 11020 26314
rect 10968 26250 11020 26256
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10140 25832 10192 25838
rect 10140 25774 10192 25780
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9496 25220 9548 25226
rect 9496 25162 9548 25168
rect 9220 24336 9272 24342
rect 9220 24278 9272 24284
rect 9508 24274 9536 25162
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9496 24268 9548 24274
rect 9496 24210 9548 24216
rect 9508 23798 9536 24210
rect 8944 23792 8996 23798
rect 8944 23734 8996 23740
rect 9496 23792 9548 23798
rect 9496 23734 9548 23740
rect 8944 23656 8996 23662
rect 8944 23598 8996 23604
rect 8956 22778 8984 23598
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9678 22944 9734 22953
rect 9508 22778 9536 22918
rect 8944 22772 8996 22778
rect 8944 22714 8996 22720
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9036 22432 9088 22438
rect 8956 22392 9036 22420
rect 8956 21554 8984 22392
rect 9036 22374 9088 22380
rect 9494 22400 9550 22409
rect 9494 22335 9550 22344
rect 9508 22234 9536 22335
rect 9600 22273 9628 22918
rect 9678 22879 9734 22888
rect 9586 22264 9642 22273
rect 9496 22228 9548 22234
rect 9586 22199 9642 22208
rect 9496 22170 9548 22176
rect 9692 22166 9720 22879
rect 9876 22817 9904 25094
rect 9968 24818 9996 25230
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 9862 22808 9918 22817
rect 9862 22743 9918 22752
rect 9864 22704 9916 22710
rect 9864 22646 9916 22652
rect 9772 22500 9824 22506
rect 9772 22442 9824 22448
rect 9784 22166 9812 22442
rect 9128 22160 9180 22166
rect 9128 22102 9180 22108
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8956 20806 8984 20946
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8482 19952 8538 19961
rect 8482 19887 8538 19896
rect 8312 18698 8432 18714
rect 8300 18692 8432 18698
rect 8352 18686 8432 18692
rect 8300 18634 8352 18640
rect 8496 17882 8524 19887
rect 8574 19544 8630 19553
rect 8574 19479 8576 19488
rect 8628 19479 8630 19488
rect 8576 19450 8628 19456
rect 8574 19272 8630 19281
rect 8574 19207 8630 19216
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8588 15706 8616 19207
rect 8680 18154 8708 19994
rect 9048 19990 9076 21422
rect 9140 21146 9168 22102
rect 9220 22024 9272 22030
rect 9496 22024 9548 22030
rect 9220 21966 9272 21972
rect 9494 21992 9496 22001
rect 9548 21992 9550 22001
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 9140 20466 9168 21082
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9232 19990 9260 21966
rect 9494 21927 9550 21936
rect 9770 21992 9826 22001
rect 9770 21927 9772 21936
rect 9824 21927 9826 21936
rect 9772 21898 9824 21904
rect 9312 21888 9364 21894
rect 9404 21888 9456 21894
rect 9312 21830 9364 21836
rect 9402 21856 9404 21865
rect 9456 21856 9458 21865
rect 9036 19984 9088 19990
rect 9036 19926 9088 19932
rect 9220 19984 9272 19990
rect 9220 19926 9272 19932
rect 9048 19718 9076 19926
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9036 19712 9088 19718
rect 9140 19689 9168 19790
rect 9036 19654 9088 19660
rect 9126 19680 9182 19689
rect 9126 19615 9182 19624
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8772 19242 8800 19450
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 9324 19174 9352 21830
rect 9402 21791 9458 21800
rect 9586 21720 9642 21729
rect 9586 21655 9642 21664
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 9416 21078 9444 21422
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 9496 21004 9548 21010
rect 9496 20946 9548 20952
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 9416 20777 9444 20810
rect 9402 20768 9458 20777
rect 9402 20703 9458 20712
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9416 19378 9444 20198
rect 9508 20097 9536 20946
rect 9494 20088 9550 20097
rect 9494 20023 9550 20032
rect 9600 19446 9628 21655
rect 9678 21584 9734 21593
rect 9678 21519 9734 21528
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9310 18320 9366 18329
rect 8852 18284 8904 18290
rect 9310 18255 9366 18264
rect 8852 18226 8904 18232
rect 8760 18216 8812 18222
rect 8864 18193 8892 18226
rect 9324 18222 9352 18255
rect 9312 18216 9364 18222
rect 8760 18158 8812 18164
rect 8850 18184 8906 18193
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 14464 8340 14894
rect 8588 14482 8616 15438
rect 8576 14476 8628 14482
rect 8312 14436 8432 14464
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8128 13025 8156 13398
rect 8114 13016 8170 13025
rect 8114 12951 8170 12960
rect 8312 12866 8340 14282
rect 8128 12838 8340 12866
rect 8128 12209 8156 12838
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8114 12200 8170 12209
rect 8114 12135 8170 12144
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 8036 10282 8064 12038
rect 7852 10254 8064 10282
rect 7852 9926 7880 10254
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7748 8424 7800 8430
rect 7654 8392 7710 8401
rect 7748 8366 7800 8372
rect 7654 8327 7710 8336
rect 7668 6662 7696 8327
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7760 6390 7788 8366
rect 7852 6458 7880 9862
rect 7930 9072 7986 9081
rect 7930 9007 7986 9016
rect 7944 8974 7972 9007
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7944 6458 7972 8910
rect 8128 7546 8156 12135
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8220 6662 8248 12718
rect 8404 12594 8432 14436
rect 8576 14418 8628 14424
rect 8680 13394 8708 15506
rect 8772 14346 8800 18158
rect 9312 18158 9364 18164
rect 8850 18119 8906 18128
rect 9600 17678 9628 18702
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 8864 17105 8892 17614
rect 9692 17610 9720 21519
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9784 19281 9812 20402
rect 9876 20058 9904 22646
rect 9968 20942 9996 24754
rect 10048 24676 10100 24682
rect 10048 24618 10100 24624
rect 10060 24070 10088 24618
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 10060 23866 10088 24006
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 10152 22137 10180 25774
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10520 24886 10548 25638
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10508 24880 10560 24886
rect 10508 24822 10560 24828
rect 10612 24750 10640 25094
rect 10600 24744 10652 24750
rect 10600 24686 10652 24692
rect 10414 24304 10470 24313
rect 10414 24239 10470 24248
rect 10322 24032 10378 24041
rect 10322 23967 10378 23976
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10244 22642 10272 23054
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10336 22574 10364 23967
rect 10428 23662 10456 24239
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 10508 23588 10560 23594
rect 10508 23530 10560 23536
rect 10416 23248 10468 23254
rect 10414 23216 10416 23225
rect 10468 23216 10470 23225
rect 10414 23151 10470 23160
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10138 22128 10194 22137
rect 10138 22063 10194 22072
rect 10416 22024 10468 22030
rect 10152 21984 10416 22012
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9968 19854 9996 20878
rect 10060 20466 10088 21830
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 10048 20256 10100 20262
rect 10046 20224 10048 20233
rect 10100 20224 10102 20233
rect 10046 20159 10102 20168
rect 10152 20058 10180 21984
rect 10416 21966 10468 21972
rect 10416 21616 10468 21622
rect 10416 21558 10468 21564
rect 10428 20602 10456 21558
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9770 19272 9826 19281
rect 9770 19207 9826 19216
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 8850 17096 8906 17105
rect 8850 17031 8906 17040
rect 8864 16590 8892 17031
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8864 13530 8892 16526
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8680 12617 8708 12650
rect 8666 12608 8722 12617
rect 8404 12566 8616 12594
rect 8404 12170 8432 12566
rect 8482 12472 8538 12481
rect 8482 12407 8538 12416
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 8298 11928 8354 11937
rect 8298 11863 8354 11872
rect 8312 11830 8340 11863
rect 8300 11824 8352 11830
rect 8496 11778 8524 12407
rect 8300 11766 8352 11772
rect 8404 11750 8524 11778
rect 8404 11082 8432 11750
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8312 10266 8340 10542
rect 8496 10266 8524 10678
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8390 9752 8446 9761
rect 8390 9687 8392 9696
rect 8444 9687 8446 9696
rect 8392 9658 8444 9664
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 7886 8340 9318
rect 8496 9178 8524 9930
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8404 8673 8432 8978
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8390 8664 8446 8673
rect 8390 8599 8446 8608
rect 8496 8498 8524 8910
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8496 7886 8524 8434
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7760 5846 7788 6326
rect 8496 6186 8524 7822
rect 8588 6866 8616 12566
rect 8666 12543 8722 12552
rect 8956 12481 8984 15642
rect 8942 12472 8998 12481
rect 8942 12407 8998 12416
rect 8666 12336 8722 12345
rect 8666 12271 8668 12280
rect 8720 12271 8722 12280
rect 8668 12242 8720 12248
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8680 9654 8708 12106
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8680 7002 8708 9590
rect 8772 9586 8800 12174
rect 9048 11082 9076 16186
rect 9232 13530 9260 17206
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9140 13258 9168 13466
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8772 8974 8800 9522
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8864 9178 8892 9386
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7750 8984 7822
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 9048 6458 9076 11018
rect 9140 9722 9168 13194
rect 9324 12442 9352 16118
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9416 14618 9444 14894
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9508 14385 9536 15370
rect 9494 14376 9550 14385
rect 9494 14311 9550 14320
rect 9588 14272 9640 14278
rect 9416 14232 9588 14260
rect 9416 13802 9444 14232
rect 9588 14214 9640 14220
rect 9494 14104 9550 14113
rect 9494 14039 9550 14048
rect 9508 13802 9536 14039
rect 9784 14006 9812 18294
rect 9876 18290 9904 18770
rect 9968 18766 9996 19790
rect 10152 19334 10180 19994
rect 10060 19306 10180 19334
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 10060 17542 10088 19306
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10152 18426 10180 18566
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10244 17338 10272 20538
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10336 17184 10364 20402
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10428 19378 10456 19722
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10428 18698 10456 19110
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10428 17678 10456 18226
rect 10520 17746 10548 23530
rect 10612 23322 10640 24686
rect 10600 23316 10652 23322
rect 10600 23258 10652 23264
rect 10612 23186 10640 23258
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10704 23118 10732 25910
rect 12084 25906 12112 26862
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 12084 25809 12112 25842
rect 12070 25800 12126 25809
rect 11336 25764 11388 25770
rect 12070 25735 12126 25744
rect 11336 25706 11388 25712
rect 11244 25696 11296 25702
rect 11244 25638 11296 25644
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 10980 24954 11008 25298
rect 11256 25226 11284 25638
rect 11348 25362 11376 25706
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12176 25362 12204 25638
rect 11336 25356 11388 25362
rect 11336 25298 11388 25304
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 11244 25220 11296 25226
rect 11244 25162 11296 25168
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 11348 24750 11376 25298
rect 12268 25226 12296 26318
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 12256 25220 12308 25226
rect 12256 25162 12308 25168
rect 11624 24886 11652 25162
rect 11978 24984 12034 24993
rect 11978 24919 12034 24928
rect 11612 24880 11664 24886
rect 11612 24822 11664 24828
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10784 24132 10836 24138
rect 10784 24074 10836 24080
rect 10692 23112 10744 23118
rect 10690 23080 10692 23089
rect 10744 23080 10746 23089
rect 10690 23015 10746 23024
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10612 22506 10640 22578
rect 10600 22500 10652 22506
rect 10600 22442 10652 22448
rect 10612 21554 10640 22442
rect 10796 22098 10824 24074
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10888 23322 10916 24006
rect 11072 23798 11100 24210
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 10968 23792 11020 23798
rect 10968 23734 11020 23740
rect 11060 23792 11112 23798
rect 11060 23734 11112 23740
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10690 21992 10746 22001
rect 10888 21962 10916 22510
rect 10690 21927 10746 21936
rect 10876 21956 10928 21962
rect 10704 21622 10732 21927
rect 10876 21898 10928 21904
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10888 21554 10916 21898
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10612 20466 10640 21490
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10612 17678 10640 18702
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10428 17338 10456 17614
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10416 17196 10468 17202
rect 10336 17156 10416 17184
rect 10416 17138 10468 17144
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 14226 10088 15302
rect 10140 14272 10192 14278
rect 9876 14198 10088 14226
rect 10138 14240 10140 14249
rect 10192 14240 10194 14249
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9508 12986 9536 13738
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9232 11014 9260 11562
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10674 9260 10950
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9232 8514 9260 9998
rect 9324 8634 9352 12038
rect 9416 9518 9444 12854
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9508 12238 9536 12718
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9494 11248 9550 11257
rect 9494 11183 9496 11192
rect 9548 11183 9550 11192
rect 9496 11154 9548 11160
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9600 9722 9628 10542
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9494 9344 9550 9353
rect 9494 9279 9550 9288
rect 9508 9110 9536 9279
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9232 8498 9444 8514
rect 9232 8492 9456 8498
rect 9232 8486 9404 8492
rect 9404 8434 9456 8440
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9232 7410 9260 7822
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 9324 4622 9352 8366
rect 9416 7342 9444 8434
rect 9600 7478 9628 9658
rect 9692 9518 9720 13942
rect 9876 12442 9904 14198
rect 10138 14175 10194 14184
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9968 13326 9996 13874
rect 9956 13320 10008 13326
rect 10008 13268 10180 13274
rect 9956 13262 10180 13268
rect 9968 13246 10180 13262
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9968 12986 9996 13126
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9862 12336 9918 12345
rect 9862 12271 9864 12280
rect 9916 12271 9918 12280
rect 9864 12242 9916 12248
rect 9968 12238 9996 12786
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9784 9994 9812 12174
rect 10152 11914 10180 13246
rect 10244 12050 10272 16118
rect 10322 16008 10378 16017
rect 10322 15943 10324 15952
rect 10376 15943 10378 15952
rect 10324 15914 10376 15920
rect 10428 15858 10456 17138
rect 10336 15830 10456 15858
rect 10336 15162 10364 15830
rect 10612 15586 10640 17614
rect 10704 16998 10732 20402
rect 10796 17882 10824 20470
rect 10888 19854 10916 21490
rect 10980 21146 11008 23734
rect 11072 22710 11100 23734
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11244 23248 11296 23254
rect 11244 23190 11296 23196
rect 11256 23050 11284 23190
rect 11244 23044 11296 23050
rect 11244 22986 11296 22992
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 10968 21140 11020 21146
rect 10968 21082 11020 21088
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10980 19666 11008 20810
rect 11072 19825 11100 22374
rect 11164 22234 11192 22374
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11164 21078 11192 21558
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 11256 20942 11284 21966
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11256 20806 11284 20878
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11058 19816 11114 19825
rect 11058 19751 11114 19760
rect 10888 19638 11008 19666
rect 10888 18290 10916 19638
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10888 17814 10916 18226
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16182 10732 16934
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10796 16114 10824 16390
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10888 15706 10916 17750
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 10966 16144 11022 16153
rect 10966 16079 10968 16088
rect 11020 16079 11022 16088
rect 10968 16050 11020 16056
rect 10980 15881 11008 16050
rect 10966 15872 11022 15881
rect 10966 15807 11022 15816
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10428 15558 10640 15586
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10336 13818 10364 15098
rect 10428 15026 10456 15558
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10428 13938 10456 14962
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10336 13790 10456 13818
rect 10428 13326 10456 13790
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12434 10456 13262
rect 10520 12986 10548 15438
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 15314 11100 15370
rect 10980 15286 11100 15314
rect 10980 15178 11008 15286
rect 10888 15150 11008 15178
rect 11060 15156 11112 15162
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10704 14362 10732 14894
rect 10784 14408 10836 14414
rect 10704 14356 10784 14362
rect 10704 14350 10836 14356
rect 10704 14334 10824 14350
rect 10598 13832 10654 13841
rect 10598 13767 10654 13776
rect 10612 13734 10640 13767
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10428 12406 10640 12434
rect 10244 12022 10548 12050
rect 10048 11892 10100 11898
rect 10152 11886 10364 11914
rect 10048 11834 10100 11840
rect 10060 11801 10088 11834
rect 10336 11830 10364 11886
rect 10324 11824 10376 11830
rect 10046 11792 10102 11801
rect 10324 11766 10376 11772
rect 10046 11727 10102 11736
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9680 8968 9732 8974
rect 9784 8956 9812 9930
rect 9876 9654 9904 11018
rect 10244 10538 10272 11698
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 9042 9904 9318
rect 10060 9110 10088 9454
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9732 8928 9812 8956
rect 10140 8968 10192 8974
rect 9680 8910 9732 8916
rect 10140 8910 10192 8916
rect 9692 8566 9720 8910
rect 10152 8566 10180 8910
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9416 6730 9444 7278
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9692 6458 9720 7210
rect 9784 7206 9812 7346
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9784 5778 9812 7142
rect 10244 6866 10272 10474
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9602 10456 9998
rect 10336 9586 10456 9602
rect 10324 9580 10456 9586
rect 10376 9574 10456 9580
rect 10324 9522 10376 9528
rect 10336 7206 10364 9522
rect 10520 9450 10548 12022
rect 10612 10996 10640 12406
rect 10704 12238 10732 14334
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 13977 10824 14214
rect 10782 13968 10838 13977
rect 10782 13903 10838 13912
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11370 10732 12174
rect 10796 11558 10824 13903
rect 10888 13841 10916 15150
rect 11060 15098 11112 15104
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10874 13832 10930 13841
rect 10874 13767 10930 13776
rect 10980 12442 11008 15030
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10704 11342 10824 11370
rect 10692 11008 10744 11014
rect 10612 10968 10692 10996
rect 10612 10130 10640 10968
rect 10692 10950 10744 10956
rect 10796 10198 10824 11342
rect 10888 10674 10916 11766
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10612 9926 10640 10066
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10612 8974 10640 9862
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10428 7546 10456 8502
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10612 7274 10640 8910
rect 10980 8090 11008 12038
rect 11072 9178 11100 15098
rect 11164 13734 11192 17138
rect 11256 16454 11284 20742
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11256 15026 11284 16390
rect 11348 15094 11376 23598
rect 11612 23248 11664 23254
rect 11440 23196 11612 23202
rect 11440 23190 11664 23196
rect 11440 23174 11652 23190
rect 11440 23050 11468 23174
rect 11428 23044 11480 23050
rect 11428 22986 11480 22992
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 11440 19922 11468 22986
rect 11532 22234 11560 22986
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11518 21992 11574 22001
rect 11518 21927 11574 21936
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11440 19378 11468 19858
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11532 17377 11560 21927
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11518 17368 11574 17377
rect 11624 17338 11652 17546
rect 11518 17303 11574 17312
rect 11612 17332 11664 17338
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11348 14958 11376 15030
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13394 11192 13670
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11532 13326 11560 17303
rect 11612 17274 11664 17280
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11348 8634 11376 13262
rect 11716 12306 11744 23598
rect 11808 23594 11836 23802
rect 11796 23588 11848 23594
rect 11796 23530 11848 23536
rect 11900 21690 11928 24822
rect 11992 23225 12020 24919
rect 12164 24268 12216 24274
rect 12164 24210 12216 24216
rect 11978 23216 12034 23225
rect 11978 23151 12034 23160
rect 11992 22642 12020 23151
rect 12176 23050 12204 24210
rect 12268 23254 12296 25162
rect 12348 24676 12400 24682
rect 12348 24618 12400 24624
rect 12360 23662 12388 24618
rect 12452 24274 12480 26454
rect 12636 26382 12664 27542
rect 12912 26450 12940 31282
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 13188 30394 13216 30670
rect 13176 30388 13228 30394
rect 13176 30330 13228 30336
rect 13832 27062 13860 32778
rect 13912 28552 13964 28558
rect 13912 28494 13964 28500
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 12900 26444 12952 26450
rect 12900 26386 12952 26392
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12912 26234 12940 26386
rect 12728 26206 12940 26234
rect 12728 25838 12756 26206
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 12716 25832 12768 25838
rect 12716 25774 12768 25780
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12348 23656 12400 23662
rect 12440 23656 12492 23662
rect 12400 23604 12440 23610
rect 12348 23598 12492 23604
rect 12360 23582 12480 23598
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 12348 23248 12400 23254
rect 12348 23190 12400 23196
rect 12164 23044 12216 23050
rect 12164 22986 12216 22992
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 11796 20392 11848 20398
rect 11796 20334 11848 20340
rect 11808 19922 11836 20334
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 11808 18834 11836 19858
rect 11900 19786 11928 20742
rect 11992 19990 12020 21966
rect 12176 20040 12204 22986
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 12268 21146 12296 22646
rect 12360 22438 12388 23190
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12544 21672 12572 25434
rect 12728 24342 12756 25774
rect 13280 24750 13308 25910
rect 13360 25832 13412 25838
rect 13360 25774 13412 25780
rect 13372 25430 13400 25774
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13360 25424 13412 25430
rect 13360 25366 13412 25372
rect 13636 25288 13688 25294
rect 13636 25230 13688 25236
rect 13544 24880 13596 24886
rect 13544 24822 13596 24828
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 13004 24342 13032 24550
rect 12716 24336 12768 24342
rect 12716 24278 12768 24284
rect 12992 24336 13044 24342
rect 12992 24278 13044 24284
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12636 21690 12664 24006
rect 12820 23798 12848 24210
rect 12808 23792 12860 23798
rect 12808 23734 12860 23740
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13096 23610 13124 23666
rect 12820 23582 13124 23610
rect 12452 21644 12572 21672
rect 12624 21684 12676 21690
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12360 20466 12388 21354
rect 12452 21010 12480 21644
rect 12624 21626 12676 21632
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12452 20534 12480 20946
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12176 20012 12296 20040
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 12084 19378 12112 19722
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11886 19272 11942 19281
rect 11886 19207 11888 19216
rect 11940 19207 11942 19216
rect 11888 19178 11940 19184
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11900 18034 11928 19178
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12084 18358 12112 19110
rect 12176 18698 12204 19858
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 12176 18204 12204 18634
rect 12084 18176 12204 18204
rect 11808 18006 11928 18034
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11808 15026 11836 18006
rect 11992 17270 12020 18022
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11900 15162 11928 17206
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11808 14822 11836 14962
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 12084 14346 12112 18176
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12176 17134 12204 17682
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12176 15473 12204 17070
rect 12162 15464 12218 15473
rect 12162 15399 12218 15408
rect 12176 15366 12204 15399
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 11992 14074 12020 14282
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12084 12306 12112 14282
rect 12268 13870 12296 20012
rect 12360 14482 12388 20402
rect 12544 20398 12572 21490
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 20806 12756 21286
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12636 19446 12664 20198
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12728 19310 12756 20198
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12452 19122 12480 19178
rect 12452 19094 12572 19122
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12452 17542 12480 18158
rect 12544 17882 12572 19094
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 18358 12664 18566
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12728 17678 12756 19246
rect 12820 19242 12848 23582
rect 13188 22506 13216 24210
rect 13372 23168 13400 24686
rect 13556 24410 13584 24822
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13280 23140 13400 23168
rect 13452 23180 13504 23186
rect 13176 22500 13228 22506
rect 13176 22442 13228 22448
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12912 20534 12940 21830
rect 12992 21004 13044 21010
rect 12992 20946 13044 20952
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12544 16658 12572 16730
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12544 14618 12572 14826
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11440 11830 11468 12106
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11624 10606 11652 12242
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11716 11540 11744 11698
rect 11808 11694 11836 12038
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11716 11512 11836 11540
rect 11808 11150 11836 11512
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11624 8430 11652 10542
rect 11716 8634 11744 10678
rect 11808 9994 11836 11086
rect 12176 10962 12204 13194
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12084 10934 12204 10962
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11900 10130 11928 10202
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11900 8566 11928 10066
rect 11992 9994 12020 10406
rect 12084 10130 12112 10934
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 12084 9654 12112 10066
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10612 6866 10640 7210
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 11900 6730 11928 8502
rect 11992 8344 12020 9522
rect 12360 8956 12388 13126
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12544 11286 12572 11630
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12636 11014 12664 17546
rect 13004 17218 13032 20946
rect 13096 20874 13124 22374
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13096 18698 13124 19654
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 13188 18222 13216 22442
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13280 17746 13308 23140
rect 13452 23122 13504 23128
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 13372 22710 13400 22986
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 13360 22500 13412 22506
rect 13360 22442 13412 22448
rect 13372 21010 13400 22442
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13358 20904 13414 20913
rect 13358 20839 13414 20848
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 12912 17190 13032 17218
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15434 12848 15846
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12820 12986 12848 13942
rect 12912 13802 12940 17190
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 13004 16046 13032 17070
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 13096 15434 13124 17546
rect 13280 17066 13308 17682
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 14618 13032 15302
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12912 12986 12940 13738
rect 13188 13258 13216 16594
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13280 14890 13308 15098
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 13004 12170 13032 12650
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 13188 11898 13216 12854
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 12714 11384 12770 11393
rect 12714 11319 12716 11328
rect 12768 11319 12770 11328
rect 12716 11290 12768 11296
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12728 10538 12756 11086
rect 13280 10674 13308 14826
rect 13372 14414 13400 20839
rect 13464 20398 13492 23122
rect 13544 23044 13596 23050
rect 13544 22986 13596 22992
rect 13556 22234 13584 22986
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13648 22098 13676 25230
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 13740 22642 13768 24278
rect 13832 24070 13860 25638
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13728 22636 13780 22642
rect 13728 22578 13780 22584
rect 13740 22506 13768 22578
rect 13728 22500 13780 22506
rect 13728 22442 13780 22448
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13648 20942 13676 21558
rect 13740 21486 13768 22034
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13636 20936 13688 20942
rect 13636 20878 13688 20884
rect 13740 20602 13768 21422
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13464 19922 13492 20334
rect 13832 20058 13860 23802
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13452 19916 13504 19922
rect 13504 19876 13584 19904
rect 13452 19858 13504 19864
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13464 19514 13492 19722
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13556 19378 13584 19876
rect 13728 19780 13780 19786
rect 13648 19740 13728 19768
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13648 19258 13676 19740
rect 13728 19722 13780 19728
rect 13464 19230 13676 19258
rect 13464 15162 13492 19230
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13556 14414 13584 18838
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13648 17270 13676 18158
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 13740 16250 13768 18294
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13648 14618 13676 15030
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13372 13954 13400 14350
rect 13372 13926 13492 13954
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13372 12714 13400 13806
rect 13464 13326 13492 13926
rect 13556 13462 13584 14350
rect 13636 14272 13688 14278
rect 13634 14240 13636 14249
rect 13688 14240 13690 14249
rect 13634 14175 13690 14184
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13188 9994 13216 10406
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 13004 9450 13032 9658
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12452 8956 12480 9046
rect 12360 8945 12480 8956
rect 12346 8936 12480 8945
rect 12402 8928 12480 8936
rect 12716 8968 12768 8974
rect 12346 8871 12402 8880
rect 12544 8916 12716 8922
rect 12544 8910 12768 8916
rect 12544 8894 12756 8910
rect 12544 8838 12572 8894
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12452 8401 12480 8570
rect 12438 8392 12494 8401
rect 11992 8316 12296 8344
rect 12438 8327 12494 8336
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7852 2446 7880 2790
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 9232 2378 9260 4422
rect 11992 2582 12020 7686
rect 12268 7546 12296 8316
rect 13096 8022 13124 9522
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12268 5642 12296 7482
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 13004 2650 13032 7346
rect 13188 6730 13216 9318
rect 13464 8634 13492 13262
rect 13648 12442 13676 14175
rect 13832 13326 13860 14826
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13740 12714 13768 13194
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13740 8090 13768 10610
rect 13832 10130 13860 11290
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13820 9580 13872 9586
rect 13924 9568 13952 28494
rect 14016 21570 14044 36518
rect 14464 27328 14516 27334
rect 14464 27270 14516 27276
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14924 27328 14976 27334
rect 14924 27270 14976 27276
rect 14188 27056 14240 27062
rect 14188 26998 14240 27004
rect 14096 25220 14148 25226
rect 14096 25162 14148 25168
rect 14108 24138 14136 25162
rect 14200 24818 14228 26998
rect 14372 26240 14424 26246
rect 14372 26182 14424 26188
rect 14384 25974 14412 26182
rect 14372 25968 14424 25974
rect 14372 25910 14424 25916
rect 14476 25226 14504 27270
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14464 25220 14516 25226
rect 14464 25162 14516 25168
rect 14476 25129 14504 25162
rect 14462 25120 14518 25129
rect 14462 25055 14518 25064
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14200 24274 14228 24754
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 14476 24138 14504 24618
rect 14096 24132 14148 24138
rect 14096 24074 14148 24080
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14108 23866 14136 24074
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14108 22030 14136 23802
rect 14292 23254 14320 23285
rect 14280 23248 14332 23254
rect 14568 23202 14596 26318
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 14752 24750 14780 25434
rect 14844 25294 14872 27270
rect 14936 27062 14964 27270
rect 14924 27056 14976 27062
rect 14924 26998 14976 27004
rect 15028 26042 15056 37062
rect 16132 29306 16160 37266
rect 16776 37126 16804 39200
rect 18064 37262 18092 39200
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 18880 37256 18932 37262
rect 18880 37198 18932 37204
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 16120 29300 16172 29306
rect 16120 29242 16172 29248
rect 15660 29028 15712 29034
rect 15660 28970 15712 28976
rect 15568 27940 15620 27946
rect 15568 27882 15620 27888
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15488 27470 15516 27814
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 15304 25838 15332 26318
rect 15384 26308 15436 26314
rect 15384 26250 15436 26256
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 14832 25288 14884 25294
rect 14832 25230 14884 25236
rect 14844 24993 14872 25230
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15304 24993 15332 25094
rect 14830 24984 14886 24993
rect 14830 24919 14886 24928
rect 15290 24984 15346 24993
rect 15396 24954 15424 26250
rect 15488 25226 15516 27406
rect 15580 25906 15608 27882
rect 15672 27062 15700 28970
rect 16868 28762 16896 37198
rect 18144 37120 18196 37126
rect 18144 37062 18196 37068
rect 18156 36786 18184 37062
rect 18144 36780 18196 36786
rect 18144 36722 18196 36728
rect 17684 36372 17736 36378
rect 17684 36314 17736 36320
rect 17696 35894 17724 36314
rect 17328 35866 17724 35894
rect 17224 29504 17276 29510
rect 17224 29446 17276 29452
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16396 27396 16448 27402
rect 16396 27338 16448 27344
rect 15660 27056 15712 27062
rect 15660 26998 15712 27004
rect 16408 26994 16436 27338
rect 16672 27056 16724 27062
rect 16672 26998 16724 27004
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 15844 26920 15896 26926
rect 15844 26862 15896 26868
rect 15856 26450 15884 26862
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15476 25220 15528 25226
rect 15476 25162 15528 25168
rect 15290 24919 15346 24928
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14752 24426 14780 24686
rect 14332 23196 14596 23202
rect 14280 23190 14596 23196
rect 14292 23174 14596 23190
rect 14660 24398 14780 24426
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14188 21616 14240 21622
rect 14016 21542 14136 21570
rect 14188 21558 14240 21564
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 14016 19310 14044 21354
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14108 18902 14136 21542
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 14016 12782 14044 18634
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14108 16046 14136 17070
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14200 15570 14228 21558
rect 14292 21486 14320 23174
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 14292 19922 14320 20266
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14292 18766 14320 19858
rect 14384 19718 14412 23054
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22710 14504 22918
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14476 21622 14504 22034
rect 14464 21616 14516 21622
rect 14464 21558 14516 21564
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14476 20890 14504 21422
rect 14660 21418 14688 24398
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14752 23118 14780 24278
rect 14844 23526 14872 24822
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14556 20936 14608 20942
rect 14476 20884 14556 20890
rect 14476 20878 14608 20884
rect 14476 20862 14596 20878
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14384 18426 14412 18906
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14292 16522 14320 16934
rect 14280 16516 14332 16522
rect 14280 16458 14332 16464
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14016 12102 14044 12310
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13872 9540 13952 9568
rect 13820 9522 13872 9528
rect 14016 9217 14044 11698
rect 14108 10742 14136 15438
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14200 13870 14228 14894
rect 14384 14074 14412 16118
rect 14476 15706 14504 19790
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14660 16590 14688 19314
rect 14752 19310 14780 23054
rect 14936 22574 14964 23598
rect 15108 23180 15160 23186
rect 15108 23122 15160 23128
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 14936 22438 14964 22510
rect 15120 22506 15148 23122
rect 15108 22500 15160 22506
rect 15108 22442 15160 22448
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 14936 22098 14964 22170
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 15120 21622 15148 22442
rect 15198 22128 15254 22137
rect 15198 22063 15200 22072
rect 15252 22063 15254 22072
rect 15200 22034 15252 22040
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 15016 21412 15068 21418
rect 15016 21354 15068 21360
rect 15028 21146 15056 21354
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 14936 20262 14964 20538
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14844 17610 14872 19382
rect 15028 19378 15056 21082
rect 15212 20602 15240 21898
rect 15396 21622 15424 24890
rect 15488 24018 15516 25162
rect 15580 24410 15608 25842
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15488 23990 15700 24018
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15488 22234 15516 22374
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15384 21072 15436 21078
rect 15384 21014 15436 21020
rect 15396 20874 15424 21014
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15120 20058 15148 20470
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14936 17490 14964 19246
rect 14844 17462 14964 17490
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14476 15586 14504 15642
rect 14476 15558 14596 15586
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14476 14414 14504 14894
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14108 9926 14136 10678
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14002 9208 14058 9217
rect 14002 9143 14058 9152
rect 14016 8634 14044 9143
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 14108 7954 14136 9862
rect 14200 8022 14228 13806
rect 14292 13530 14320 13942
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14292 11354 14320 12718
rect 14384 12442 14412 12854
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14464 12232 14516 12238
rect 14462 12200 14464 12209
rect 14516 12200 14518 12209
rect 14462 12135 14518 12144
rect 14568 11762 14596 15558
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14476 11642 14504 11698
rect 14476 11614 14596 11642
rect 14568 11558 14596 11614
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14476 11082 14504 11494
rect 14660 11234 14688 16390
rect 14844 14006 14872 17462
rect 15028 16998 15056 19314
rect 15212 18834 15240 19654
rect 15304 18970 15332 20402
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15212 18358 15240 18770
rect 15396 18698 15424 19110
rect 15488 18834 15516 22170
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15580 20874 15608 21830
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15672 20602 15700 23990
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15856 19174 15884 26386
rect 16408 26234 16436 26930
rect 16580 26784 16632 26790
rect 16580 26726 16632 26732
rect 16408 26206 16528 26234
rect 16212 25764 16264 25770
rect 16212 25706 16264 25712
rect 16224 25498 16252 25706
rect 16212 25492 16264 25498
rect 16212 25434 16264 25440
rect 16500 25294 16528 26206
rect 16592 25838 16620 26726
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16028 25152 16080 25158
rect 16028 25094 16080 25100
rect 16040 24954 16068 25094
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 16488 24268 16540 24274
rect 16488 24210 16540 24216
rect 15936 24132 15988 24138
rect 15936 24074 15988 24080
rect 15948 23798 15976 24074
rect 16120 24064 16172 24070
rect 16120 24006 16172 24012
rect 16132 23798 16160 24006
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 15948 22098 15976 23734
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16224 22778 16252 23598
rect 16500 23118 16528 24210
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16592 23186 16620 24074
rect 16684 23322 16712 26998
rect 17236 26586 17264 29446
rect 17224 26580 17276 26586
rect 17224 26522 17276 26528
rect 16856 26240 16908 26246
rect 16856 26182 16908 26188
rect 16948 26240 17000 26246
rect 16948 26182 17000 26188
rect 16868 23322 16896 26182
rect 16960 24177 16988 26182
rect 17040 25968 17092 25974
rect 17040 25910 17092 25916
rect 17052 25498 17080 25910
rect 17236 25838 17264 26522
rect 17328 26450 17356 35866
rect 18892 33114 18920 37198
rect 19996 37126 20024 39200
rect 21284 37126 21312 39200
rect 22008 37256 22060 37262
rect 22008 37198 22060 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 18880 33108 18932 33114
rect 18880 33050 18932 33056
rect 18236 32904 18288 32910
rect 18236 32846 18288 32852
rect 17592 26920 17644 26926
rect 17592 26862 17644 26868
rect 17500 26512 17552 26518
rect 17500 26454 17552 26460
rect 17316 26444 17368 26450
rect 17316 26386 17368 26392
rect 17224 25832 17276 25838
rect 17224 25774 17276 25780
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 17132 24880 17184 24886
rect 17132 24822 17184 24828
rect 17052 24313 17080 24822
rect 17144 24750 17172 24822
rect 17328 24750 17356 26386
rect 17512 26228 17540 26454
rect 17604 26314 17632 26862
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17420 26200 17540 26228
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17038 24304 17094 24313
rect 17038 24239 17094 24248
rect 17224 24200 17276 24206
rect 16946 24168 17002 24177
rect 17224 24142 17276 24148
rect 16946 24103 17002 24112
rect 17236 24041 17264 24142
rect 17222 24032 17278 24041
rect 17222 23967 17278 23976
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 15936 22092 15988 22098
rect 16500 22094 16528 23054
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 15936 22034 15988 22040
rect 16040 22066 16528 22094
rect 16040 20448 16068 22066
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16224 21622 16252 21966
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 15948 20420 16068 20448
rect 15948 19530 15976 20420
rect 16026 20360 16082 20369
rect 16026 20295 16028 20304
rect 16080 20295 16082 20304
rect 16028 20266 16080 20272
rect 15948 19502 16068 19530
rect 16132 19514 16160 21558
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 16394 21040 16450 21049
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 15212 17746 15240 18294
rect 15304 18222 15332 18566
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14936 13258 14964 15982
rect 15120 15162 15148 17070
rect 15304 16046 15332 18158
rect 15948 17542 15976 19314
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 15396 16250 15424 17206
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 15028 14618 15056 15030
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 15120 13870 15148 15098
rect 15304 14618 15332 15370
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 15120 12434 15148 13806
rect 15304 13462 15332 14214
rect 15396 13530 15424 15030
rect 15580 14006 15608 15506
rect 15672 14958 15700 16594
rect 15856 16522 15884 16934
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15488 13530 15516 13942
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15028 12406 15148 12434
rect 14922 12200 14978 12209
rect 14922 12135 14978 12144
rect 14568 11206 14688 11234
rect 14832 11212 14884 11218
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14568 10810 14596 11206
rect 14832 11154 14884 11160
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14292 9994 14320 10474
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9450 14320 9930
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14568 8634 14596 9522
rect 14660 9518 14688 11018
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14752 9042 14780 10678
rect 14844 10470 14872 11154
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14844 9178 14872 9930
rect 14936 9178 14964 12135
rect 15028 9654 15056 12406
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15212 10062 15240 11698
rect 15396 11218 15424 12582
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15488 11898 15516 12106
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15474 11792 15530 11801
rect 15474 11727 15476 11736
rect 15528 11727 15530 11736
rect 15476 11698 15528 11704
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 15120 8838 15148 9522
rect 15488 9382 15516 11698
rect 15580 11014 15608 12106
rect 15672 12102 15700 14894
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15672 10606 15700 12038
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15764 10538 15792 15370
rect 15948 12442 15976 17478
rect 16040 15910 16068 19502
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16132 19242 16160 19314
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16132 14618 16160 16050
rect 16224 16046 16252 21014
rect 16394 20975 16450 20984
rect 16488 21004 16540 21010
rect 16408 20942 16436 20975
rect 16488 20946 16540 20952
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16316 15570 16344 20742
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16408 17746 16436 19314
rect 16500 18902 16528 20946
rect 16776 20534 16804 22374
rect 17052 21690 17080 23734
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17236 21962 17264 23598
rect 17328 23118 17356 24550
rect 17420 23798 17448 26200
rect 17512 26042 17540 26200
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17500 25832 17552 25838
rect 17500 25774 17552 25780
rect 17512 24274 17540 25774
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17408 23792 17460 23798
rect 17408 23734 17460 23740
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16868 21350 16896 21490
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16856 20936 16908 20942
rect 16854 20904 16856 20913
rect 16908 20904 16910 20913
rect 16854 20839 16910 20848
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16592 19718 16620 20402
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 18970 16620 19654
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16776 18290 16804 20470
rect 17144 20058 17172 21898
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16776 17814 16804 18226
rect 16764 17808 16816 17814
rect 16764 17750 16816 17756
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16408 17270 16436 17682
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15948 12102 15976 12378
rect 16132 12345 16160 14554
rect 16408 14414 16436 17002
rect 16868 16114 16896 19994
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16960 18834 16988 19246
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16960 16250 16988 16458
rect 17236 16250 17264 20198
rect 17328 19990 17356 23054
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 17512 17270 17540 23462
rect 17604 22094 17632 26250
rect 18248 25906 18276 32846
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 17776 25696 17828 25702
rect 17776 25638 17828 25644
rect 18144 25696 18196 25702
rect 18144 25638 18196 25644
rect 17788 25226 17816 25638
rect 17868 25424 17920 25430
rect 17868 25366 17920 25372
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 17880 25106 17908 25366
rect 18156 25362 18184 25638
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 18052 25152 18104 25158
rect 17788 25078 17908 25106
rect 17972 25112 18052 25140
rect 17788 24886 17816 25078
rect 17776 24880 17828 24886
rect 17776 24822 17828 24828
rect 17788 23254 17816 24822
rect 17972 24138 18000 25112
rect 18052 25094 18104 25100
rect 18156 24274 18184 25298
rect 18524 24818 18552 26250
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 18800 24818 18828 25094
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 17776 23248 17828 23254
rect 17776 23190 17828 23196
rect 17604 22066 17724 22094
rect 17592 21344 17644 21350
rect 17592 21286 17644 21292
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16118 12336 16174 12345
rect 16118 12271 16174 12280
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16224 11898 16252 12718
rect 16592 12714 16620 15914
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16776 15094 16804 15302
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 17236 14958 17264 16186
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17328 15706 17356 16118
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17236 13410 17264 14894
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 17144 13382 17264 13410
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16592 12306 16620 12650
rect 16684 12442 16712 12854
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15856 10266 15884 10678
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13280 6458 13308 6666
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 3252 800 3280 2246
rect 4540 800 4568 2246
rect 6472 800 6500 2246
rect 7760 800 7788 2246
rect 9692 800 9720 2314
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 1986 11100 2246
rect 10980 1958 11100 1986
rect 10980 800 11008 1958
rect 12912 800 12940 2382
rect 14200 800 14228 2382
rect 15120 2310 15148 8774
rect 15948 3534 15976 11154
rect 16500 9926 16528 11698
rect 16592 11218 16620 12242
rect 16776 12238 16804 13330
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11694 16804 12174
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16868 11558 16896 12378
rect 17144 11830 17172 13382
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17236 12782 17264 13194
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17328 12594 17356 15438
rect 17512 15008 17540 15846
rect 17604 15434 17632 21286
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17592 15020 17644 15026
rect 17512 14980 17592 15008
rect 17592 14962 17644 14968
rect 17696 14804 17724 22066
rect 17788 18442 17816 23190
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17880 21350 17908 23054
rect 18064 22778 18092 24074
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 17972 21894 18000 22510
rect 18616 22166 18644 24754
rect 19260 24614 19288 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 19260 24206 19288 24550
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 18800 23730 18828 24142
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18800 22982 18828 23666
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19536 23186 19564 23598
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19628 23050 19656 23462
rect 19616 23044 19668 23050
rect 19616 22986 19668 22992
rect 18788 22976 18840 22982
rect 18786 22944 18788 22953
rect 18840 22944 18842 22953
rect 18786 22879 18842 22888
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19628 22234 19656 22374
rect 19616 22228 19668 22234
rect 19616 22170 19668 22176
rect 18052 22160 18104 22166
rect 18052 22102 18104 22108
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 18064 19334 18092 22102
rect 20088 22094 20116 25434
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20824 24410 20852 25162
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 20812 24404 20864 24410
rect 20812 24346 20864 24352
rect 21100 24070 21128 24754
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 20272 23798 20300 24006
rect 20260 23792 20312 23798
rect 20260 23734 20312 23740
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20272 22438 20300 22578
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20088 22066 20208 22094
rect 18236 21956 18288 21962
rect 18236 21898 18288 21904
rect 19248 21956 19300 21962
rect 19248 21898 19300 21904
rect 18248 21146 18276 21898
rect 18788 21412 18840 21418
rect 18788 21354 18840 21360
rect 18800 21146 18828 21354
rect 18236 21140 18288 21146
rect 18236 21082 18288 21088
rect 18788 21140 18840 21146
rect 18788 21082 18840 21088
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18432 19854 18460 20198
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18156 19446 18184 19654
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18432 19378 18460 19790
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18420 19372 18472 19378
rect 18064 19306 18184 19334
rect 18420 19314 18472 19320
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17788 18414 17908 18442
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17512 14776 17724 14804
rect 17408 13864 17460 13870
rect 17512 13852 17540 14776
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17460 13824 17540 13852
rect 17408 13806 17460 13812
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17420 12986 17448 13194
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17236 12566 17356 12594
rect 17236 12209 17264 12566
rect 17420 12374 17448 12922
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17222 12200 17278 12209
rect 17222 12135 17278 12144
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 17420 11393 17448 11766
rect 17406 11384 17462 11393
rect 17512 11354 17540 13824
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17604 11830 17632 12038
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17406 11319 17462 11328
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9722 16528 9862
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16868 8906 16896 11018
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16960 8634 16988 10542
rect 17052 9926 17080 11222
rect 17512 11082 17540 11290
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17604 11014 17632 11630
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10674 17632 10950
rect 17696 10810 17724 13874
rect 17788 12170 17816 15302
rect 17880 15162 17908 18414
rect 17972 18086 18000 18634
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 13938 17908 14214
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17972 13530 18000 15030
rect 18064 14482 18092 16662
rect 18156 15609 18184 19306
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18248 16590 18276 17546
rect 18432 17066 18460 19314
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18340 16658 18368 16934
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 15910 18552 16526
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18142 15600 18198 15609
rect 18142 15535 18198 15544
rect 18156 15502 18184 15535
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18616 15094 18644 19722
rect 18800 19446 18828 21082
rect 19260 20874 19288 21898
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 19076 19378 19104 19926
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18788 18692 18840 18698
rect 18788 18634 18840 18640
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 18708 15706 18736 18634
rect 18800 18426 18828 18634
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18880 17060 18932 17066
rect 18880 17002 18932 17008
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18800 15434 18828 15846
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18052 14476 18104 14482
rect 18104 14436 18276 14464
rect 18052 14418 18104 14424
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 17776 12164 17828 12170
rect 17776 12106 17828 12112
rect 17868 11620 17920 11626
rect 17868 11562 17920 11568
rect 17880 11286 17908 11562
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 18064 11082 18092 11494
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 18156 10130 18184 12718
rect 18248 11694 18276 14436
rect 18340 12850 18368 14962
rect 18418 13968 18474 13977
rect 18418 13903 18420 13912
rect 18472 13903 18474 13912
rect 18420 13874 18472 13880
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18524 10742 18552 11494
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6458 17264 6598
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17696 5370 17724 9658
rect 18616 9518 18644 15030
rect 18800 14618 18828 15370
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18800 13938 18828 14554
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18800 13530 18828 13874
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18800 12646 18828 13262
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 17512 2446 17540 4966
rect 18616 3058 18644 8434
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18616 2650 18644 2994
rect 18892 2990 18920 17002
rect 18984 16794 19012 18634
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 19076 17542 19104 18226
rect 19260 18222 19288 20810
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 19514 19380 20742
rect 19444 19990 19472 21422
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19628 19786 19656 20266
rect 20180 19786 20208 22066
rect 20272 20466 20300 22374
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20732 21894 20760 21966
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20272 20058 20300 20402
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19720 18714 19748 19314
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19720 18686 19840 18714
rect 19812 18630 19840 18686
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19352 17762 19380 18022
rect 19444 17882 19472 18294
rect 19996 18086 20024 19246
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 20180 18222 20208 18770
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19352 17734 19472 17762
rect 19444 17678 19472 17734
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18970 15600 19026 15609
rect 18970 15535 19026 15544
rect 18984 15502 19012 15535
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18984 13462 19012 13670
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 12442 19012 12582
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 19076 2582 19104 17478
rect 19444 16998 19472 17614
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19628 16658 19656 17070
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19720 16726 19748 16934
rect 19812 16794 19840 16934
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19708 16720 19760 16726
rect 19708 16662 19760 16668
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19352 16182 19380 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19800 16176 19852 16182
rect 19800 16118 19852 16124
rect 19812 15502 19840 16118
rect 19904 15638 19932 16186
rect 19892 15632 19944 15638
rect 19892 15574 19944 15580
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 14482 20024 18022
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 20180 17542 20208 17750
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 20088 14958 20116 15982
rect 20180 15978 20208 17478
rect 20352 16720 20404 16726
rect 20352 16662 20404 16668
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 20076 14340 20128 14346
rect 20076 14282 20128 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19248 13796 19300 13802
rect 19248 13738 19300 13744
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19168 12918 19196 13670
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19260 12782 19288 13738
rect 19996 13326 20024 13942
rect 20088 13530 20116 14282
rect 20180 13870 20208 15914
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20272 15094 20300 15506
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19444 11898 19472 12854
rect 19996 12850 20024 13262
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20088 12170 20116 12582
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 20272 11830 20300 12854
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19352 6798 19380 11018
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 19444 2446 19472 10406
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 20364 3466 20392 16662
rect 20456 15586 20484 19858
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20548 17746 20576 19722
rect 20628 18896 20680 18902
rect 20628 18838 20680 18844
rect 20640 18698 20668 18838
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20548 16250 20576 16526
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20640 16046 20668 18158
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20640 15638 20668 15982
rect 20628 15632 20680 15638
rect 20456 15558 20576 15586
rect 20628 15574 20680 15580
rect 20444 15428 20496 15434
rect 20444 15370 20496 15376
rect 20456 15162 20484 15370
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20548 12918 20576 15558
rect 20732 15026 20760 21830
rect 21100 19310 21128 24006
rect 21192 22710 21220 30670
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 21180 22704 21232 22710
rect 21180 22646 21232 22652
rect 21284 21894 21312 23598
rect 22020 21962 22048 37198
rect 23216 37126 23244 39200
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 22560 30048 22612 30054
rect 22560 29990 22612 29996
rect 22572 26450 22600 29990
rect 22560 26444 22612 26450
rect 22560 26386 22612 26392
rect 22572 25362 22600 26386
rect 22560 25356 22612 25362
rect 22560 25298 22612 25304
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21824 21888 21876 21894
rect 21824 21830 21876 21836
rect 21836 20874 21864 21830
rect 21916 21412 21968 21418
rect 21916 21354 21968 21360
rect 21824 20868 21876 20874
rect 21824 20810 21876 20816
rect 21272 19440 21324 19446
rect 21272 19382 21324 19388
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21100 18290 21128 19246
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 21008 17490 21036 17546
rect 21008 17462 21128 17490
rect 21100 17270 21128 17462
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 21008 16794 21036 17206
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14482 20668 14894
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20536 12912 20588 12918
rect 20536 12854 20588 12860
rect 20824 11898 20852 13398
rect 20916 13394 20944 15438
rect 21192 15094 21220 18634
rect 21284 18426 21312 19382
rect 21836 18834 21864 20810
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21732 18148 21784 18154
rect 21732 18090 21784 18096
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21652 17338 21680 17682
rect 21640 17332 21692 17338
rect 21640 17274 21692 17280
rect 21744 17134 21772 18090
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21468 16794 21496 17002
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16794 21588 16934
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21284 14822 21312 14962
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21744 14346 21772 17070
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21008 13462 21036 13874
rect 20996 13456 21048 13462
rect 20996 13398 21048 13404
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 21100 12102 21128 14282
rect 21652 13530 21680 14282
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 21836 10810 21864 17614
rect 21928 16726 21956 21354
rect 23308 20602 23336 37198
rect 24504 37126 24532 39200
rect 26436 37466 26464 39200
rect 26424 37460 26476 37466
rect 26424 37402 26476 37408
rect 26424 37324 26476 37330
rect 26424 37266 26476 37272
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 24596 30938 24624 37198
rect 26436 36174 26464 37266
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 27448 36854 27476 37198
rect 27724 37126 27752 39200
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 29092 37256 29144 37262
rect 29092 37198 29144 37204
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 28460 36922 28488 37198
rect 29104 36922 29132 37198
rect 29656 37126 29684 39200
rect 30944 37126 30972 39200
rect 32876 37466 32904 39200
rect 34164 37466 34192 39200
rect 35530 38176 35586 38185
rect 35530 38111 35586 38120
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 32864 37460 32916 37466
rect 32864 37402 32916 37408
rect 34152 37460 34204 37466
rect 34152 37402 34204 37408
rect 32956 37324 33008 37330
rect 32956 37266 33008 37272
rect 34796 37324 34848 37330
rect 34796 37266 34848 37272
rect 31024 37256 31076 37262
rect 31024 37198 31076 37204
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 30932 37120 30984 37126
rect 30932 37062 30984 37068
rect 28448 36916 28500 36922
rect 28448 36858 28500 36864
rect 29092 36916 29144 36922
rect 29092 36858 29144 36864
rect 27436 36848 27488 36854
rect 27436 36790 27488 36796
rect 27160 36780 27212 36786
rect 27160 36722 27212 36728
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 27172 35086 27200 36722
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 27172 29646 27200 35022
rect 27448 30258 27476 36790
rect 28356 36576 28408 36582
rect 28356 36518 28408 36524
rect 28368 36378 28396 36518
rect 28356 36372 28408 36378
rect 28356 36314 28408 36320
rect 31036 32842 31064 37198
rect 31024 32836 31076 32842
rect 31024 32778 31076 32784
rect 27804 31816 27856 31822
rect 27804 31758 27856 31764
rect 27436 30252 27488 30258
rect 27436 30194 27488 30200
rect 27160 29640 27212 29646
rect 27160 29582 27212 29588
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23768 23118 23796 23462
rect 24688 23322 24716 24074
rect 27816 23866 27844 31758
rect 32968 30122 32996 37266
rect 32956 30116 33008 30122
rect 32956 30058 33008 30064
rect 33784 24948 33836 24954
rect 33784 24890 33836 24896
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 24676 23316 24728 23322
rect 24676 23258 24728 23264
rect 24688 23118 24716 23258
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 22466 19952 22522 19961
rect 22466 19887 22522 19896
rect 22480 19854 22508 19887
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22204 19446 22232 19654
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22112 17882 22140 19246
rect 22940 18426 22968 19790
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 22940 18290 22968 18362
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21916 16720 21968 16726
rect 21916 16662 21968 16668
rect 22112 14006 22140 17818
rect 22388 17814 22416 18022
rect 22376 17808 22428 17814
rect 22376 17750 22428 17756
rect 22480 16998 22508 18226
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22558 16144 22614 16153
rect 22558 16079 22560 16088
rect 22612 16079 22614 16088
rect 22560 16050 22612 16056
rect 22572 15706 22600 16050
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22190 15464 22246 15473
rect 22190 15399 22192 15408
rect 22244 15399 22246 15408
rect 22192 15370 22244 15376
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22204 13326 22232 14486
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22480 14074 22508 14282
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22756 13938 22784 14214
rect 23492 14006 23520 14758
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22480 13530 22508 13806
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 23400 13326 23428 13874
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 22204 12986 22232 13262
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22100 12708 22152 12714
rect 22100 12650 22152 12656
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 22112 6322 22140 12650
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20640 2514 20668 2790
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 20732 2446 20760 3334
rect 23676 2582 23704 22918
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24872 18902 24900 22578
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 27632 18358 27660 23666
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27160 9376 27212 9382
rect 27160 9318 27212 9324
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24584 6180 24636 6186
rect 24584 6122 24636 6128
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 24596 2446 24624 6122
rect 24688 2446 24716 6598
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 25700 2378 25728 4082
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 27080 2378 27108 2790
rect 27172 2582 27200 9318
rect 29840 2650 29868 18906
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 29828 2644 29880 2650
rect 29828 2586 29880 2592
rect 27160 2576 27212 2582
rect 27160 2518 27212 2524
rect 30392 2446 30420 2790
rect 30576 2650 30604 15642
rect 32404 14000 32456 14006
rect 32404 13942 32456 13948
rect 32416 2650 32444 13942
rect 33796 2650 33824 24890
rect 34808 24138 34836 37266
rect 35544 36922 35572 38111
rect 35624 37256 35676 37262
rect 35624 37198 35676 37204
rect 35532 36916 35584 36922
rect 35532 36858 35584 36864
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35636 36378 35664 37198
rect 36096 37126 36124 39200
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 37384 36854 37412 39200
rect 37372 36848 37424 36854
rect 37372 36790 37424 36796
rect 36176 36576 36228 36582
rect 36176 36518 36228 36524
rect 35624 36372 35676 36378
rect 35624 36314 35676 36320
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35636 26234 35664 36314
rect 36188 35894 36216 36518
rect 36266 36136 36322 36145
rect 36266 36071 36322 36080
rect 36280 36038 36308 36071
rect 36268 36032 36320 36038
rect 36268 35974 36320 35980
rect 36188 35866 36492 35894
rect 36360 35080 36412 35086
rect 36360 35022 36412 35028
rect 36372 34785 36400 35022
rect 36358 34776 36414 34785
rect 36358 34711 36360 34720
rect 36412 34711 36414 34720
rect 36360 34682 36412 34688
rect 36268 32836 36320 32842
rect 36268 32778 36320 32784
rect 36280 32745 36308 32778
rect 36266 32736 36322 32745
rect 36266 32671 36322 32680
rect 35808 31952 35860 31958
rect 35808 31894 35860 31900
rect 35820 31385 35848 31894
rect 35806 31376 35862 31385
rect 35806 31311 35862 31320
rect 36268 29572 36320 29578
rect 36268 29514 36320 29520
rect 35992 29504 36044 29510
rect 35992 29446 36044 29452
rect 35900 27940 35952 27946
rect 35900 27882 35952 27888
rect 35808 26512 35860 26518
rect 35808 26454 35860 26460
rect 35544 26206 35664 26234
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 24132 34848 24138
rect 34796 24074 34848 24080
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34520 20256 34572 20262
rect 34520 20198 34572 20204
rect 34532 18290 34560 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34520 18284 34572 18290
rect 34520 18226 34572 18232
rect 30564 2644 30616 2650
rect 30564 2586 30616 2592
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 33784 2644 33836 2650
rect 33784 2586 33836 2592
rect 34532 2582 34560 18226
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35544 16017 35572 26206
rect 35820 25945 35848 26454
rect 35806 25936 35862 25945
rect 35912 25906 35940 27882
rect 35806 25871 35862 25880
rect 35900 25900 35952 25906
rect 35900 25842 35952 25848
rect 35900 24744 35952 24750
rect 35900 24686 35952 24692
rect 35912 22030 35940 24686
rect 35900 22024 35952 22030
rect 35900 21966 35952 21972
rect 35912 19378 35940 21966
rect 36004 21418 36032 29446
rect 36280 29345 36308 29514
rect 36266 29336 36322 29345
rect 36266 29271 36322 29280
rect 36268 28076 36320 28082
rect 36268 28018 36320 28024
rect 36280 27985 36308 28018
rect 36266 27976 36322 27985
rect 36266 27911 36322 27920
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 35992 21412 36044 21418
rect 35992 21354 36044 21360
rect 36096 20602 36124 26318
rect 36360 24744 36412 24750
rect 36360 24686 36412 24692
rect 36372 24585 36400 24686
rect 36358 24576 36414 24585
rect 36358 24511 36414 24520
rect 36372 24410 36400 24511
rect 36360 24404 36412 24410
rect 36360 24346 36412 24352
rect 36266 22536 36322 22545
rect 36266 22471 36268 22480
rect 36320 22471 36322 22480
rect 36268 22442 36320 22448
rect 36268 21548 36320 21554
rect 36268 21490 36320 21496
rect 36176 21344 36228 21350
rect 36176 21286 36228 21292
rect 36188 20806 36216 21286
rect 36280 21185 36308 21490
rect 36266 21176 36322 21185
rect 36266 21111 36322 21120
rect 36176 20800 36228 20806
rect 36176 20742 36228 20748
rect 36084 20596 36136 20602
rect 36084 20538 36136 20544
rect 35900 19372 35952 19378
rect 35900 19314 35952 19320
rect 36084 19168 36136 19174
rect 36084 19110 36136 19116
rect 36096 18290 36124 19110
rect 36084 18284 36136 18290
rect 36084 18226 36136 18232
rect 36268 18080 36320 18086
rect 36268 18022 36320 18028
rect 36280 17785 36308 18022
rect 36266 17776 36322 17785
rect 36266 17711 36322 17720
rect 36464 16726 36492 35866
rect 36544 32768 36596 32774
rect 36544 32710 36596 32716
rect 36556 17542 36584 32710
rect 36636 20052 36688 20058
rect 36636 19994 36688 20000
rect 36544 17536 36596 17542
rect 36544 17478 36596 17484
rect 36452 16720 36504 16726
rect 36452 16662 36504 16668
rect 36360 16108 36412 16114
rect 36360 16050 36412 16056
rect 35530 16008 35586 16017
rect 35530 15943 35586 15952
rect 35900 15904 35952 15910
rect 35900 15846 35952 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35532 14272 35584 14278
rect 35532 14214 35584 14220
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35544 12306 35572 14214
rect 35912 13326 35940 15846
rect 36372 15745 36400 16050
rect 36358 15736 36414 15745
rect 36358 15671 36414 15680
rect 36266 14376 36322 14385
rect 36266 14311 36322 14320
rect 36280 14278 36308 14311
rect 36268 14272 36320 14278
rect 36268 14214 36320 14220
rect 35900 13320 35952 13326
rect 35900 13262 35952 13268
rect 36084 13184 36136 13190
rect 36084 13126 36136 13132
rect 35808 12844 35860 12850
rect 35808 12786 35860 12792
rect 35820 12345 35848 12786
rect 35806 12336 35862 12345
rect 35532 12300 35584 12306
rect 35806 12271 35862 12280
rect 35532 12242 35584 12248
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 36096 11150 36124 13126
rect 36268 11280 36320 11286
rect 36268 11222 36320 11228
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 36280 10985 36308 11222
rect 36266 10976 36322 10985
rect 36266 10911 36322 10920
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35452 3194 35480 9862
rect 36084 9716 36136 9722
rect 36084 9658 36136 9664
rect 36096 9110 36124 9658
rect 36084 9104 36136 9110
rect 36084 9046 36136 9052
rect 36266 8936 36322 8945
rect 36266 8871 36268 8880
rect 36320 8871 36322 8880
rect 36268 8842 36320 8848
rect 36648 8090 36676 19994
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36268 7812 36320 7818
rect 36268 7754 36320 7760
rect 36280 7585 36308 7754
rect 36266 7576 36322 7585
rect 36266 7511 36322 7520
rect 36176 6452 36228 6458
rect 36176 6394 36228 6400
rect 35530 5672 35586 5681
rect 35530 5607 35532 5616
rect 35584 5607 35586 5616
rect 35532 5578 35584 5584
rect 36084 4616 36136 4622
rect 36084 4558 36136 4564
rect 36096 3942 36124 4558
rect 36084 3936 36136 3942
rect 36084 3878 36136 3884
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35440 3188 35492 3194
rect 35440 3130 35492 3136
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34520 2576 34572 2582
rect 34520 2518 34572 2524
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 25688 2372 25740 2378
rect 25688 2314 25740 2320
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 16132 800 16160 2314
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 17420 800 17448 2246
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20640 800 20668 2246
rect 22572 800 22600 2246
rect 23860 800 23888 2246
rect 25792 800 25820 2246
rect 27080 800 27108 2314
rect 29000 2304 29052 2310
rect 30392 2292 30420 2382
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 33508 2372 33560 2378
rect 33508 2314 33560 2320
rect 29000 2246 29052 2252
rect 30300 2264 30420 2292
rect 29012 800 29040 2246
rect 30300 800 30328 2264
rect 32232 800 32260 2314
rect 33520 800 33548 2314
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 35452 800 35480 2246
rect 35820 2145 35848 3470
rect 36188 3194 36216 6394
rect 36268 5568 36320 5574
rect 36266 5536 36268 5545
rect 36320 5536 36322 5545
rect 36266 5471 36322 5480
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 36280 4185 36308 4422
rect 36266 4176 36322 4185
rect 36266 4111 36322 4120
rect 36176 3188 36228 3194
rect 36176 3130 36228 3136
rect 36728 3120 36780 3126
rect 36728 3062 36780 3068
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 36372 2310 36400 2994
rect 36360 2304 36412 2310
rect 36360 2246 36412 2252
rect 35806 2136 35862 2145
rect 35806 2071 35862 2080
rect 36372 1465 36400 2246
rect 36358 1456 36414 1465
rect 36358 1391 36414 1400
rect 36740 800 36768 3062
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 7746 200 7802 800
rect 9678 200 9734 800
rect 10966 200 11022 800
rect 12898 200 12954 800
rect 14186 200 14242 800
rect 16118 200 16174 800
rect 17406 200 17462 800
rect 19338 200 19394 800
rect 20626 200 20682 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 33506 200 33562 800
rect 35438 200 35494 800
rect 36726 200 36782 800
<< via2 >>
rect 1674 37440 1730 37496
rect 2870 38800 2926 38856
rect 1858 36216 1914 36272
rect 1582 35400 1638 35456
rect 1582 32020 1638 32056
rect 1582 32000 1584 32020
rect 1584 32000 1636 32020
rect 1636 32000 1638 32020
rect 1674 30640 1730 30696
rect 1582 28600 1638 28656
rect 1674 27276 1676 27296
rect 1676 27276 1728 27296
rect 1728 27276 1730 27296
rect 1674 27240 1730 27276
rect 1582 23840 1638 23896
rect 1858 27412 1860 27432
rect 1860 27412 1912 27432
rect 1912 27412 1914 27432
rect 1858 27376 1914 27412
rect 1674 21836 1676 21856
rect 1676 21836 1728 21856
rect 1728 21836 1730 21856
rect 1674 21800 1730 21836
rect 1674 20440 1730 20496
rect 1674 18400 1730 18456
rect 2502 22072 2558 22128
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 3146 25200 3202 25256
rect 2778 23432 2834 23488
rect 2686 19780 2742 19816
rect 2686 19760 2688 19780
rect 2688 19760 2740 19780
rect 2740 19760 2742 19780
rect 3054 19488 3110 19544
rect 2410 17060 2466 17096
rect 2410 17040 2412 17060
rect 2412 17040 2464 17060
rect 2464 17040 2466 17060
rect 1582 9560 1638 9616
rect 2778 13640 2834 13696
rect 2870 13232 2926 13288
rect 2686 11736 2742 11792
rect 1950 8744 2006 8800
rect 1674 4800 1730 4856
rect 2318 5636 2374 5672
rect 2318 5616 2320 5636
rect 2320 5616 2372 5636
rect 2372 5616 2374 5636
rect 1674 3440 1730 3496
rect 2778 6840 2834 6896
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3790 21664 3846 21720
rect 3422 20596 3478 20632
rect 3422 20576 3424 20596
rect 3424 20576 3476 20596
rect 3476 20576 3478 20596
rect 3514 18128 3570 18184
rect 3330 12960 3386 13016
rect 3882 20576 3938 20632
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4526 19252 4528 19272
rect 4528 19252 4580 19272
rect 4580 19252 4582 19272
rect 4526 19216 4582 19252
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4710 20168 4766 20224
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 5170 20848 5226 20904
rect 5170 18828 5226 18864
rect 5170 18808 5172 18828
rect 5172 18808 5224 18828
rect 5224 18808 5226 18828
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4250 16652 4306 16688
rect 4250 16632 4252 16652
rect 4252 16632 4304 16652
rect 4304 16632 4306 16652
rect 4710 16496 4766 16552
rect 4710 16224 4766 16280
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4066 15020 4122 15056
rect 4066 15000 4068 15020
rect 4068 15000 4120 15020
rect 4120 15000 4122 15020
rect 3790 11600 3846 11656
rect 3974 10260 4030 10296
rect 3974 10240 3976 10260
rect 3976 10240 4028 10260
rect 4028 10240 4030 10260
rect 3974 8200 4030 8256
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4986 16496 5042 16552
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4894 8492 4950 8528
rect 4894 8472 4896 8492
rect 4896 8472 4948 8492
rect 4948 8472 4950 8492
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5262 18264 5318 18320
rect 5630 18944 5686 19000
rect 5446 18264 5502 18320
rect 5262 16224 5318 16280
rect 5354 12280 5410 12336
rect 6642 20712 6698 20768
rect 6826 21800 6882 21856
rect 6826 19624 6882 19680
rect 6734 18944 6790 19000
rect 5998 17040 6054 17096
rect 5998 16632 6054 16688
rect 7838 24148 7840 24168
rect 7840 24148 7892 24168
rect 7892 24148 7894 24168
rect 7838 24112 7894 24148
rect 7746 23180 7802 23216
rect 7746 23160 7748 23180
rect 7748 23160 7800 23180
rect 7800 23160 7802 23180
rect 7562 21664 7618 21720
rect 7654 21120 7710 21176
rect 7102 18808 7158 18864
rect 7470 20032 7526 20088
rect 8022 22344 8078 22400
rect 8390 22616 8446 22672
rect 8114 21120 8170 21176
rect 8022 19896 8078 19952
rect 8022 19352 8078 19408
rect 6734 15816 6790 15872
rect 6458 13388 6514 13424
rect 6458 13368 6460 13388
rect 6460 13368 6512 13388
rect 6512 13368 6514 13388
rect 6090 8900 6146 8936
rect 6090 8880 6092 8900
rect 6092 8880 6144 8900
rect 6144 8880 6146 8900
rect 6366 11192 6422 11248
rect 6642 13096 6698 13152
rect 6550 12588 6552 12608
rect 6552 12588 6604 12608
rect 6604 12588 6606 12608
rect 6550 12552 6606 12588
rect 6550 12280 6606 12336
rect 7838 17312 7894 17368
rect 6918 13368 6974 13424
rect 6734 12688 6790 12744
rect 7470 13232 7526 13288
rect 7102 13096 7158 13152
rect 7562 11892 7618 11928
rect 7562 11872 7564 11892
rect 7564 11872 7616 11892
rect 7616 11872 7618 11892
rect 7286 9696 7342 9752
rect 7194 9288 7250 9344
rect 7102 8472 7158 8528
rect 7470 9152 7526 9208
rect 7378 8744 7434 8800
rect 7470 8608 7526 8664
rect 7102 8236 7104 8256
rect 7104 8236 7156 8256
rect 7156 8236 7158 8256
rect 7102 8200 7158 8236
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 7470 6860 7526 6896
rect 7470 6840 7472 6860
rect 7472 6840 7524 6860
rect 7524 6840 7526 6860
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8574 21936 8630 21992
rect 8666 20868 8722 20904
rect 8666 20848 8668 20868
rect 8668 20848 8720 20868
rect 8720 20848 8722 20868
rect 12530 29452 12532 29472
rect 12532 29452 12584 29472
rect 12584 29452 12586 29472
rect 12530 29416 12586 29452
rect 9494 22344 9550 22400
rect 9678 22888 9734 22944
rect 9586 22208 9642 22264
rect 9862 22752 9918 22808
rect 8482 19896 8538 19952
rect 8574 19508 8630 19544
rect 8574 19488 8576 19508
rect 8576 19488 8628 19508
rect 8628 19488 8630 19508
rect 8574 19216 8630 19272
rect 9494 21972 9496 21992
rect 9496 21972 9548 21992
rect 9548 21972 9550 21992
rect 9494 21936 9550 21972
rect 9770 21956 9826 21992
rect 9770 21936 9772 21956
rect 9772 21936 9824 21956
rect 9824 21936 9826 21956
rect 9402 21836 9404 21856
rect 9404 21836 9456 21856
rect 9456 21836 9458 21856
rect 9126 19624 9182 19680
rect 9402 21800 9458 21836
rect 9586 21664 9642 21720
rect 9402 20712 9458 20768
rect 9494 20032 9550 20088
rect 9678 21528 9734 21584
rect 9310 18264 9366 18320
rect 8114 12960 8170 13016
rect 8114 12144 8170 12200
rect 7654 8336 7710 8392
rect 7930 9016 7986 9072
rect 8850 18128 8906 18184
rect 10414 24248 10470 24304
rect 10322 23976 10378 24032
rect 10414 23196 10416 23216
rect 10416 23196 10468 23216
rect 10468 23196 10470 23216
rect 10414 23160 10470 23196
rect 10138 22072 10194 22128
rect 10046 20204 10048 20224
rect 10048 20204 10100 20224
rect 10100 20204 10102 20224
rect 10046 20168 10102 20204
rect 9770 19216 9826 19272
rect 8850 17040 8906 17096
rect 8482 12416 8538 12472
rect 8298 11872 8354 11928
rect 8390 9716 8446 9752
rect 8390 9696 8392 9716
rect 8392 9696 8444 9716
rect 8444 9696 8446 9716
rect 8390 8608 8446 8664
rect 8666 12552 8722 12608
rect 8942 12416 8998 12472
rect 8666 12300 8722 12336
rect 8666 12280 8668 12300
rect 8668 12280 8720 12300
rect 8720 12280 8722 12300
rect 9494 14320 9550 14376
rect 9494 14048 9550 14104
rect 12070 25744 12126 25800
rect 11978 24928 12034 24984
rect 10690 23060 10692 23080
rect 10692 23060 10744 23080
rect 10744 23060 10746 23080
rect 10690 23024 10746 23060
rect 10690 21936 10746 21992
rect 10138 14220 10140 14240
rect 10140 14220 10192 14240
rect 10192 14220 10194 14240
rect 9494 11212 9550 11248
rect 9494 11192 9496 11212
rect 9496 11192 9548 11212
rect 9548 11192 9550 11212
rect 9494 9288 9550 9344
rect 10138 14184 10194 14220
rect 9862 12300 9918 12336
rect 9862 12280 9864 12300
rect 9864 12280 9916 12300
rect 9916 12280 9918 12300
rect 10322 15972 10378 16008
rect 10322 15952 10324 15972
rect 10324 15952 10376 15972
rect 10376 15952 10378 15972
rect 11058 19760 11114 19816
rect 10966 16108 11022 16144
rect 10966 16088 10968 16108
rect 10968 16088 11020 16108
rect 11020 16088 11022 16108
rect 10966 15816 11022 15872
rect 10598 13776 10654 13832
rect 10046 11736 10102 11792
rect 10782 13912 10838 13968
rect 10874 13776 10930 13832
rect 11518 21936 11574 21992
rect 11518 17312 11574 17368
rect 11978 23160 12034 23216
rect 11886 19236 11942 19272
rect 11886 19216 11888 19236
rect 11888 19216 11940 19236
rect 11940 19216 11942 19236
rect 12162 15408 12218 15464
rect 13358 20848 13414 20904
rect 12714 11348 12770 11384
rect 12714 11328 12716 11348
rect 12716 11328 12768 11348
rect 12768 11328 12770 11348
rect 13634 14220 13636 14240
rect 13636 14220 13688 14240
rect 13688 14220 13690 14240
rect 13634 14184 13690 14220
rect 12346 8880 12402 8936
rect 12438 8336 12494 8392
rect 14462 25064 14518 25120
rect 14830 24928 14886 24984
rect 15290 24928 15346 24984
rect 15198 22092 15254 22128
rect 15198 22072 15200 22092
rect 15200 22072 15252 22092
rect 15252 22072 15254 22092
rect 14002 9152 14058 9208
rect 14462 12180 14464 12200
rect 14464 12180 14516 12200
rect 14516 12180 14518 12200
rect 14462 12144 14518 12180
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 17038 24248 17094 24304
rect 16946 24112 17002 24168
rect 17222 23976 17278 24032
rect 16026 20324 16082 20360
rect 16026 20304 16028 20324
rect 16028 20304 16080 20324
rect 16080 20304 16082 20324
rect 14922 12144 14978 12200
rect 15474 11756 15530 11792
rect 15474 11736 15476 11756
rect 15476 11736 15528 11756
rect 15528 11736 15530 11756
rect 16394 20984 16450 21040
rect 16854 20884 16856 20904
rect 16856 20884 16908 20904
rect 16908 20884 16910 20904
rect 16854 20848 16910 20884
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 16118 12280 16174 12336
rect 1674 1400 1730 1456
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 18786 22924 18788 22944
rect 18788 22924 18840 22944
rect 18840 22924 18842 22944
rect 18786 22888 18842 22924
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 17222 12144 17278 12200
rect 17406 11328 17462 11384
rect 18142 15544 18198 15600
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 18418 13932 18474 13968
rect 18418 13912 18420 13932
rect 18420 13912 18472 13932
rect 18472 13912 18474 13932
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 18970 15544 19026 15600
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 35530 38120 35586 38176
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 22466 19896 22522 19952
rect 22558 16108 22614 16144
rect 22558 16088 22560 16108
rect 22560 16088 22612 16108
rect 22612 16088 22614 16108
rect 22190 15428 22246 15464
rect 22190 15408 22192 15428
rect 22192 15408 22244 15428
rect 22244 15408 22246 15428
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 36266 36080 36322 36136
rect 36358 34740 36414 34776
rect 36358 34720 36360 34740
rect 36360 34720 36412 34740
rect 36412 34720 36414 34740
rect 36266 32680 36322 32736
rect 35806 31320 35862 31376
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35806 25880 35862 25936
rect 36266 29280 36322 29336
rect 36266 27920 36322 27976
rect 36358 24520 36414 24576
rect 36266 22500 36322 22536
rect 36266 22480 36268 22500
rect 36268 22480 36320 22500
rect 36320 22480 36322 22500
rect 36266 21120 36322 21176
rect 36266 17720 36322 17776
rect 35530 15952 35586 16008
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 36358 15680 36414 15736
rect 36266 14320 36322 14376
rect 35806 12280 35862 12336
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 36266 10920 36322 10976
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 36266 8900 36322 8936
rect 36266 8880 36268 8900
rect 36268 8880 36320 8900
rect 36320 8880 36322 8900
rect 36266 7520 36322 7576
rect 35530 5636 35586 5672
rect 35530 5616 35532 5636
rect 35532 5616 35584 5636
rect 35584 5616 35586 5636
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 36266 5516 36268 5536
rect 36268 5516 36320 5536
rect 36320 5516 36322 5536
rect 36266 5480 36322 5516
rect 36266 4120 36322 4176
rect 35806 2080 35862 2136
rect 36358 1400 36414 1456
<< metal3 >>
rect 200 38858 800 38888
rect 2865 38858 2931 38861
rect 200 38856 2931 38858
rect 200 38800 2870 38856
rect 2926 38800 2931 38856
rect 200 38798 2931 38800
rect 200 38768 800 38798
rect 2865 38795 2931 38798
rect 35525 38178 35591 38181
rect 37200 38178 37800 38208
rect 35525 38176 37800 38178
rect 35525 38120 35530 38176
rect 35586 38120 37800 38176
rect 35525 38118 37800 38120
rect 35525 38115 35591 38118
rect 37200 38088 37800 38118
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 1669 37498 1735 37501
rect 200 37496 1735 37498
rect 200 37440 1674 37496
rect 1730 37440 1735 37496
rect 200 37438 1735 37440
rect 200 37408 800 37438
rect 1669 37435 1735 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 1853 36276 1919 36277
rect 1853 36272 1900 36276
rect 1964 36274 1970 36276
rect 1853 36216 1858 36272
rect 1853 36212 1900 36216
rect 1964 36214 2010 36274
rect 1964 36212 1970 36214
rect 1853 36211 1919 36212
rect 36261 36138 36327 36141
rect 37200 36138 37800 36168
rect 36261 36136 37800 36138
rect 36261 36080 36266 36136
rect 36322 36080 37800 36136
rect 36261 36078 37800 36080
rect 36261 36075 36327 36078
rect 37200 36048 37800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35458 800 35488
rect 1577 35458 1643 35461
rect 200 35456 1643 35458
rect 200 35400 1582 35456
rect 1638 35400 1643 35456
rect 200 35398 1643 35400
rect 200 35368 800 35398
rect 1577 35395 1643 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 36353 34778 36419 34781
rect 37200 34778 37800 34808
rect 36353 34776 37800 34778
rect 36353 34720 36358 34776
rect 36414 34720 37800 34776
rect 36353 34718 37800 34720
rect 36353 34715 36419 34718
rect 37200 34688 37800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34008 800 34128
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 36261 32738 36327 32741
rect 37200 32738 37800 32768
rect 36261 32736 37800 32738
rect 36261 32680 36266 32736
rect 36322 32680 37800 32736
rect 36261 32678 37800 32680
rect 36261 32675 36327 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 37200 32648 37800 32678
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 200 32056 1643 32058
rect 200 32000 1582 32056
rect 1638 32000 1643 32056
rect 200 31998 1643 32000
rect 200 31968 800 31998
rect 1577 31995 1643 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 35801 31378 35867 31381
rect 37200 31378 37800 31408
rect 35801 31376 37800 31378
rect 35801 31320 35806 31376
rect 35862 31320 37800 31376
rect 35801 31318 37800 31320
rect 35801 31315 35867 31318
rect 37200 31288 37800 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1669 30698 1735 30701
rect 200 30696 1735 30698
rect 200 30640 1674 30696
rect 1730 30640 1735 30696
rect 200 30638 1735 30640
rect 200 30608 800 30638
rect 1669 30635 1735 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 12525 29476 12591 29477
rect 12525 29474 12572 29476
rect 12480 29472 12572 29474
rect 12480 29416 12530 29472
rect 12480 29414 12572 29416
rect 12525 29412 12572 29414
rect 12636 29412 12642 29476
rect 12525 29411 12591 29412
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 36261 29338 36327 29341
rect 37200 29338 37800 29368
rect 36261 29336 37800 29338
rect 36261 29280 36266 29336
rect 36322 29280 37800 29336
rect 36261 29278 37800 29280
rect 36261 29275 36327 29278
rect 37200 29248 37800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1577 28658 1643 28661
rect 200 28656 1643 28658
rect 200 28600 1582 28656
rect 1638 28600 1643 28656
rect 200 28598 1643 28600
rect 200 28568 800 28598
rect 1577 28595 1643 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 36261 27978 36327 27981
rect 37200 27978 37800 28008
rect 36261 27976 37800 27978
rect 36261 27920 36266 27976
rect 36322 27920 37800 27976
rect 36261 27918 37800 27920
rect 36261 27915 36327 27918
rect 37200 27888 37800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 1853 27434 1919 27437
rect 2078 27434 2084 27436
rect 1853 27432 2084 27434
rect 1853 27376 1858 27432
rect 1914 27376 2084 27432
rect 1853 27374 2084 27376
rect 1853 27371 1919 27374
rect 2078 27372 2084 27374
rect 2148 27372 2154 27436
rect 200 27298 800 27328
rect 1669 27298 1735 27301
rect 200 27296 1735 27298
rect 200 27240 1674 27296
rect 1730 27240 1735 27296
rect 200 27238 1735 27240
rect 200 27208 800 27238
rect 1669 27235 1735 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 35801 25938 35867 25941
rect 37200 25938 37800 25968
rect 35801 25936 37800 25938
rect 35801 25880 35806 25936
rect 35862 25880 37800 25936
rect 35801 25878 37800 25880
rect 35801 25875 35867 25878
rect 37200 25848 37800 25878
rect 12065 25802 12131 25805
rect 12198 25802 12204 25804
rect 12065 25800 12204 25802
rect 12065 25744 12070 25800
rect 12126 25744 12204 25800
rect 12065 25742 12204 25744
rect 12065 25739 12131 25742
rect 12198 25740 12204 25742
rect 12268 25740 12274 25804
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 3141 25258 3207 25261
rect 200 25256 3207 25258
rect 200 25200 3146 25256
rect 3202 25200 3207 25256
rect 200 25198 3207 25200
rect 200 25168 800 25198
rect 3141 25195 3207 25198
rect 14457 25122 14523 25125
rect 14590 25122 14596 25124
rect 14457 25120 14596 25122
rect 14457 25064 14462 25120
rect 14518 25064 14596 25120
rect 14457 25062 14596 25064
rect 14457 25059 14523 25062
rect 14590 25060 14596 25062
rect 14660 25060 14666 25124
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 11973 24986 12039 24989
rect 14825 24986 14891 24989
rect 11973 24984 14891 24986
rect 11973 24928 11978 24984
rect 12034 24928 14830 24984
rect 14886 24928 14891 24984
rect 11973 24926 14891 24928
rect 11973 24923 12039 24926
rect 14825 24923 14891 24926
rect 15285 24988 15351 24989
rect 15285 24984 15332 24988
rect 15396 24986 15402 24988
rect 15285 24928 15290 24984
rect 15285 24924 15332 24928
rect 15396 24926 15442 24986
rect 15396 24924 15402 24926
rect 15285 24923 15351 24924
rect 36353 24578 36419 24581
rect 37200 24578 37800 24608
rect 36353 24576 37800 24578
rect 36353 24520 36358 24576
rect 36414 24520 37800 24576
rect 36353 24518 37800 24520
rect 36353 24515 36419 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 37200 24488 37800 24518
rect 34930 24447 35246 24448
rect 10409 24306 10475 24309
rect 17033 24306 17099 24309
rect 10409 24304 17099 24306
rect 10409 24248 10414 24304
rect 10470 24248 17038 24304
rect 17094 24248 17099 24304
rect 10409 24246 17099 24248
rect 10409 24243 10475 24246
rect 17033 24243 17099 24246
rect 7833 24170 7899 24173
rect 16941 24170 17007 24173
rect 7833 24168 17007 24170
rect 7833 24112 7838 24168
rect 7894 24112 16946 24168
rect 17002 24112 17007 24168
rect 7833 24110 17007 24112
rect 7833 24107 7899 24110
rect 16941 24107 17007 24110
rect 10317 24034 10383 24037
rect 17217 24034 17283 24037
rect 10317 24032 17283 24034
rect 10317 23976 10322 24032
rect 10378 23976 17222 24032
rect 17278 23976 17283 24032
rect 10317 23974 17283 23976
rect 10317 23971 10383 23974
rect 17217 23971 17283 23974
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1577 23898 1643 23901
rect 200 23896 1643 23898
rect 200 23840 1582 23896
rect 1638 23840 1643 23896
rect 200 23838 1643 23840
rect 200 23808 800 23838
rect 1577 23835 1643 23838
rect 2773 23492 2839 23493
rect 2773 23488 2820 23492
rect 2884 23490 2890 23492
rect 2773 23432 2778 23488
rect 2773 23428 2820 23432
rect 2884 23430 2930 23490
rect 2884 23428 2890 23430
rect 2773 23427 2839 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 1894 23156 1900 23220
rect 1964 23218 1970 23220
rect 7741 23218 7807 23221
rect 1964 23216 7807 23218
rect 1964 23160 7746 23216
rect 7802 23160 7807 23216
rect 1964 23158 7807 23160
rect 1964 23156 1970 23158
rect 7741 23155 7807 23158
rect 10409 23218 10475 23221
rect 11973 23218 12039 23221
rect 10409 23216 12039 23218
rect 10409 23160 10414 23216
rect 10470 23160 11978 23216
rect 12034 23160 12039 23216
rect 10409 23158 12039 23160
rect 10409 23155 10475 23158
rect 11973 23155 12039 23158
rect 10685 23084 10751 23085
rect 10685 23080 10732 23084
rect 10796 23082 10802 23084
rect 10685 23024 10690 23080
rect 10685 23020 10732 23024
rect 10796 23022 10842 23082
rect 10796 23020 10802 23022
rect 10685 23019 10751 23020
rect 9673 22946 9739 22949
rect 18781 22946 18847 22949
rect 9673 22944 18847 22946
rect 9673 22888 9678 22944
rect 9734 22888 18786 22944
rect 18842 22888 18847 22944
rect 9673 22886 18847 22888
rect 9673 22883 9739 22886
rect 18781 22883 18847 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 9857 22812 9923 22813
rect 9806 22810 9812 22812
rect 9766 22750 9812 22810
rect 9876 22808 9923 22812
rect 9918 22752 9923 22808
rect 9806 22748 9812 22750
rect 9876 22748 9923 22752
rect 9857 22747 9923 22748
rect 8385 22676 8451 22677
rect 8334 22674 8340 22676
rect 8294 22614 8340 22674
rect 8404 22672 8451 22676
rect 8446 22616 8451 22672
rect 8334 22612 8340 22614
rect 8404 22612 8451 22616
rect 8385 22611 8451 22612
rect 36261 22538 36327 22541
rect 37200 22538 37800 22568
rect 36261 22536 37800 22538
rect 36261 22480 36266 22536
rect 36322 22480 37800 22536
rect 36261 22478 37800 22480
rect 36261 22475 36327 22478
rect 37200 22448 37800 22478
rect 8017 22402 8083 22405
rect 9489 22402 9555 22405
rect 8017 22400 9555 22402
rect 8017 22344 8022 22400
rect 8078 22344 9494 22400
rect 9550 22344 9555 22400
rect 8017 22342 9555 22344
rect 8017 22339 8083 22342
rect 9489 22339 9555 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 9581 22266 9647 22269
rect 9581 22264 9690 22266
rect 9581 22208 9586 22264
rect 9642 22208 9690 22264
rect 9581 22203 9690 22208
rect 2497 22130 2563 22133
rect 4654 22130 4660 22132
rect 2497 22128 4660 22130
rect 2497 22072 2502 22128
rect 2558 22072 4660 22128
rect 2497 22070 4660 22072
rect 2497 22067 2563 22070
rect 4654 22068 4660 22070
rect 4724 22068 4730 22132
rect 8569 21994 8635 21997
rect 9489 21994 9555 21997
rect 8569 21992 9555 21994
rect 8569 21936 8574 21992
rect 8630 21936 9494 21992
rect 9550 21936 9555 21992
rect 8569 21934 9555 21936
rect 8569 21931 8635 21934
rect 9489 21931 9555 21934
rect 200 21858 800 21888
rect 1669 21858 1735 21861
rect 200 21856 1735 21858
rect 200 21800 1674 21856
rect 1730 21800 1735 21856
rect 200 21798 1735 21800
rect 200 21768 800 21798
rect 1669 21795 1735 21798
rect 6821 21858 6887 21861
rect 7966 21858 7972 21860
rect 6821 21856 7972 21858
rect 6821 21800 6826 21856
rect 6882 21800 7972 21856
rect 6821 21798 7972 21800
rect 6821 21795 6887 21798
rect 7966 21796 7972 21798
rect 8036 21858 8042 21860
rect 9397 21858 9463 21861
rect 8036 21856 9463 21858
rect 8036 21800 9402 21856
rect 9458 21800 9463 21856
rect 8036 21798 9463 21800
rect 8036 21796 8042 21798
rect 9397 21795 9463 21798
rect 9630 21725 9690 22203
rect 10133 22130 10199 22133
rect 15193 22130 15259 22133
rect 10133 22128 15259 22130
rect 10133 22072 10138 22128
rect 10194 22072 15198 22128
rect 15254 22072 15259 22128
rect 10133 22070 15259 22072
rect 10133 22067 10199 22070
rect 9765 21994 9831 21997
rect 10685 21994 10751 21997
rect 9765 21992 10751 21994
rect 9765 21936 9770 21992
rect 9826 21936 10690 21992
rect 10746 21936 10751 21992
rect 9765 21934 10751 21936
rect 9765 21931 9831 21934
rect 10685 21931 10751 21934
rect 11513 21994 11579 21997
rect 11654 21994 11714 22070
rect 15193 22067 15259 22070
rect 11513 21992 11714 21994
rect 11513 21936 11518 21992
rect 11574 21936 11714 21992
rect 11513 21934 11714 21936
rect 11513 21931 11579 21934
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 3785 21722 3851 21725
rect 7557 21722 7623 21725
rect 3785 21720 7623 21722
rect 3785 21664 3790 21720
rect 3846 21664 7562 21720
rect 7618 21664 7623 21720
rect 3785 21662 7623 21664
rect 3785 21659 3851 21662
rect 7557 21659 7623 21662
rect 9581 21720 9690 21725
rect 9581 21664 9586 21720
rect 9642 21664 9690 21720
rect 9581 21662 9690 21664
rect 9581 21659 9647 21662
rect 9673 21586 9739 21589
rect 9806 21586 9812 21588
rect 9673 21584 9812 21586
rect 9673 21528 9678 21584
rect 9734 21528 9812 21584
rect 9673 21526 9812 21528
rect 9673 21523 9739 21526
rect 9806 21524 9812 21526
rect 9876 21524 9882 21588
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 7649 21178 7715 21181
rect 8109 21178 8175 21181
rect 7649 21176 8175 21178
rect 7649 21120 7654 21176
rect 7710 21120 8114 21176
rect 8170 21120 8175 21176
rect 7649 21118 8175 21120
rect 7649 21115 7715 21118
rect 8109 21115 8175 21118
rect 36261 21178 36327 21181
rect 37200 21178 37800 21208
rect 36261 21176 37800 21178
rect 36261 21120 36266 21176
rect 36322 21120 37800 21176
rect 36261 21118 37800 21120
rect 36261 21115 36327 21118
rect 37200 21088 37800 21118
rect 12566 20980 12572 21044
rect 12636 21042 12642 21044
rect 16389 21042 16455 21045
rect 12636 21040 16455 21042
rect 12636 20984 16394 21040
rect 16450 20984 16455 21040
rect 12636 20982 16455 20984
rect 12636 20980 12642 20982
rect 16389 20979 16455 20982
rect 5165 20906 5231 20909
rect 8661 20908 8727 20909
rect 8661 20906 8708 20908
rect 5165 20904 8708 20906
rect 8772 20906 8778 20908
rect 13353 20906 13419 20909
rect 16849 20906 16915 20909
rect 5165 20848 5170 20904
rect 5226 20848 8666 20904
rect 5165 20846 8708 20848
rect 5165 20843 5231 20846
rect 8661 20844 8708 20846
rect 8772 20846 8854 20906
rect 13353 20904 16915 20906
rect 13353 20848 13358 20904
rect 13414 20848 16854 20904
rect 16910 20848 16915 20904
rect 13353 20846 16915 20848
rect 8772 20844 8778 20846
rect 8661 20843 8727 20844
rect 13353 20843 13419 20846
rect 16849 20843 16915 20846
rect 6637 20770 6703 20773
rect 9397 20770 9463 20773
rect 6637 20768 9463 20770
rect 6637 20712 6642 20768
rect 6698 20712 9402 20768
rect 9458 20712 9463 20768
rect 6637 20710 9463 20712
rect 6637 20707 6703 20710
rect 9397 20707 9463 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 3417 20634 3483 20637
rect 3877 20634 3943 20637
rect 8334 20634 8340 20636
rect 3417 20632 8340 20634
rect 3417 20576 3422 20632
rect 3478 20576 3882 20632
rect 3938 20576 8340 20632
rect 3417 20574 8340 20576
rect 3417 20571 3483 20574
rect 3877 20571 3943 20574
rect 8334 20572 8340 20574
rect 8404 20572 8410 20636
rect 200 20498 800 20528
rect 1669 20498 1735 20501
rect 200 20496 1735 20498
rect 200 20440 1674 20496
rect 1730 20440 1735 20496
rect 200 20438 1735 20440
rect 200 20408 800 20438
rect 1669 20435 1735 20438
rect 2078 20300 2084 20364
rect 2148 20362 2154 20364
rect 16021 20362 16087 20365
rect 2148 20360 16087 20362
rect 2148 20304 16026 20360
rect 16082 20304 16087 20360
rect 2148 20302 16087 20304
rect 2148 20300 2154 20302
rect 16021 20299 16087 20302
rect 4705 20226 4771 20229
rect 10041 20226 10107 20229
rect 4705 20224 10107 20226
rect 4705 20168 4710 20224
rect 4766 20168 10046 20224
rect 10102 20168 10107 20224
rect 4705 20166 10107 20168
rect 4705 20163 4771 20166
rect 10041 20163 10107 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 7465 20090 7531 20093
rect 9489 20090 9555 20093
rect 7465 20088 9555 20090
rect 7465 20032 7470 20088
rect 7526 20032 9494 20088
rect 9550 20032 9555 20088
rect 7465 20030 9555 20032
rect 7465 20027 7531 20030
rect 9489 20027 9555 20030
rect 8017 19954 8083 19957
rect 8477 19954 8543 19957
rect 8017 19952 8543 19954
rect 8017 19896 8022 19952
rect 8078 19896 8482 19952
rect 8538 19896 8543 19952
rect 8017 19894 8543 19896
rect 8017 19891 8083 19894
rect 8477 19891 8543 19894
rect 8702 19892 8708 19956
rect 8772 19954 8778 19956
rect 22461 19954 22527 19957
rect 8772 19952 22527 19954
rect 8772 19896 22466 19952
rect 22522 19896 22527 19952
rect 8772 19894 22527 19896
rect 8772 19892 8778 19894
rect 22461 19891 22527 19894
rect 2681 19818 2747 19821
rect 11053 19818 11119 19821
rect 2681 19816 11119 19818
rect 2681 19760 2686 19816
rect 2742 19760 11058 19816
rect 11114 19760 11119 19816
rect 2681 19758 11119 19760
rect 2681 19755 2747 19758
rect 11053 19755 11119 19758
rect 6821 19682 6887 19685
rect 9121 19682 9187 19685
rect 6821 19680 9187 19682
rect 6821 19624 6826 19680
rect 6882 19624 9126 19680
rect 9182 19624 9187 19680
rect 6821 19622 9187 19624
rect 6821 19619 6887 19622
rect 9121 19619 9187 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 3049 19546 3115 19549
rect 8569 19546 8635 19549
rect 3049 19544 8635 19546
rect 3049 19488 3054 19544
rect 3110 19488 8574 19544
rect 8630 19488 8635 19544
rect 3049 19486 8635 19488
rect 3049 19483 3115 19486
rect 8569 19483 8635 19486
rect 8017 19412 8083 19413
rect 7966 19348 7972 19412
rect 8036 19410 8083 19412
rect 8036 19408 8128 19410
rect 8078 19352 8128 19408
rect 8036 19350 8128 19352
rect 8036 19348 8083 19350
rect 8017 19347 8083 19348
rect 4521 19274 4587 19277
rect 4654 19274 4660 19276
rect 4521 19272 4660 19274
rect 4521 19216 4526 19272
rect 4582 19216 4660 19272
rect 4521 19214 4660 19216
rect 4521 19211 4587 19214
rect 4654 19212 4660 19214
rect 4724 19212 4730 19276
rect 8569 19274 8635 19277
rect 9765 19274 9831 19277
rect 8569 19272 9831 19274
rect 8569 19216 8574 19272
rect 8630 19216 9770 19272
rect 9826 19216 9831 19272
rect 8569 19214 9831 19216
rect 8569 19211 8635 19214
rect 9765 19211 9831 19214
rect 11881 19274 11947 19277
rect 12198 19274 12204 19276
rect 11881 19272 12204 19274
rect 11881 19216 11886 19272
rect 11942 19216 12204 19272
rect 11881 19214 12204 19216
rect 11881 19211 11947 19214
rect 12198 19212 12204 19214
rect 12268 19212 12274 19276
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 37200 19048 37800 19168
rect 34930 19007 35246 19008
rect 5625 19002 5691 19005
rect 6729 19002 6795 19005
rect 5625 19000 6795 19002
rect 5625 18944 5630 19000
rect 5686 18944 6734 19000
rect 6790 18944 6795 19000
rect 5625 18942 6795 18944
rect 5625 18939 5691 18942
rect 6729 18939 6795 18942
rect 5165 18866 5231 18869
rect 7097 18866 7163 18869
rect 5165 18864 7163 18866
rect 5165 18808 5170 18864
rect 5226 18808 7102 18864
rect 7158 18808 7163 18864
rect 5165 18806 7163 18808
rect 5165 18803 5231 18806
rect 7097 18803 7163 18806
rect 19570 18528 19886 18529
rect 200 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 1669 18458 1735 18461
rect 200 18456 1735 18458
rect 200 18400 1674 18456
rect 1730 18400 1735 18456
rect 200 18398 1735 18400
rect 200 18368 800 18398
rect 1669 18395 1735 18398
rect 5257 18322 5323 18325
rect 5441 18322 5507 18325
rect 9305 18322 9371 18325
rect 5257 18320 9371 18322
rect 5257 18264 5262 18320
rect 5318 18264 5446 18320
rect 5502 18264 9310 18320
rect 9366 18264 9371 18320
rect 5257 18262 9371 18264
rect 5257 18259 5323 18262
rect 5441 18259 5507 18262
rect 9305 18259 9371 18262
rect 3509 18186 3575 18189
rect 8845 18186 8911 18189
rect 3509 18184 8911 18186
rect 3509 18128 3514 18184
rect 3570 18128 8850 18184
rect 8906 18128 8911 18184
rect 3509 18126 8911 18128
rect 3509 18123 3575 18126
rect 8845 18123 8911 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 36261 17778 36327 17781
rect 37200 17778 37800 17808
rect 36261 17776 37800 17778
rect 36261 17720 36266 17776
rect 36322 17720 37800 17776
rect 36261 17718 37800 17720
rect 36261 17715 36327 17718
rect 37200 17688 37800 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 7833 17370 7899 17373
rect 11513 17370 11579 17373
rect 7833 17368 11579 17370
rect 7833 17312 7838 17368
rect 7894 17312 11518 17368
rect 11574 17312 11579 17368
rect 7833 17310 11579 17312
rect 7833 17307 7899 17310
rect 11513 17307 11579 17310
rect 200 17098 800 17128
rect 2405 17098 2471 17101
rect 200 17096 2471 17098
rect 200 17040 2410 17096
rect 2466 17040 2471 17096
rect 200 17038 2471 17040
rect 200 17008 800 17038
rect 2405 17035 2471 17038
rect 5993 17098 6059 17101
rect 8845 17098 8911 17101
rect 5993 17096 8911 17098
rect 5993 17040 5998 17096
rect 6054 17040 8850 17096
rect 8906 17040 8911 17096
rect 5993 17038 8911 17040
rect 5993 17035 6059 17038
rect 8845 17035 8911 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 4245 16690 4311 16693
rect 5993 16690 6059 16693
rect 4245 16688 6059 16690
rect 4245 16632 4250 16688
rect 4306 16632 5998 16688
rect 6054 16632 6059 16688
rect 4245 16630 6059 16632
rect 4245 16627 4311 16630
rect 5993 16627 6059 16630
rect 4705 16554 4771 16557
rect 4981 16554 5047 16557
rect 4705 16552 5047 16554
rect 4705 16496 4710 16552
rect 4766 16496 4986 16552
rect 5042 16496 5047 16552
rect 4705 16494 5047 16496
rect 4705 16491 4771 16494
rect 4981 16491 5047 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4705 16282 4771 16285
rect 5257 16282 5323 16285
rect 4705 16280 5323 16282
rect 4705 16224 4710 16280
rect 4766 16224 5262 16280
rect 5318 16224 5323 16280
rect 4705 16222 5323 16224
rect 4705 16219 4771 16222
rect 5257 16219 5323 16222
rect 10961 16146 11027 16149
rect 22553 16146 22619 16149
rect 10961 16144 22619 16146
rect 10961 16088 10966 16144
rect 11022 16088 22558 16144
rect 22614 16088 22619 16144
rect 10961 16086 22619 16088
rect 10961 16083 11027 16086
rect 22553 16083 22619 16086
rect 10317 16010 10383 16013
rect 35525 16010 35591 16013
rect 10317 16008 35591 16010
rect 10317 15952 10322 16008
rect 10378 15952 35530 16008
rect 35586 15952 35591 16008
rect 10317 15950 35591 15952
rect 10317 15947 10383 15950
rect 35525 15947 35591 15950
rect 6729 15874 6795 15877
rect 10961 15874 11027 15877
rect 6729 15872 11027 15874
rect 6729 15816 6734 15872
rect 6790 15816 10966 15872
rect 11022 15816 11027 15872
rect 6729 15814 11027 15816
rect 6729 15811 6795 15814
rect 10961 15811 11027 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 36353 15738 36419 15741
rect 37200 15738 37800 15768
rect 36353 15736 37800 15738
rect 36353 15680 36358 15736
rect 36414 15680 37800 15736
rect 36353 15678 37800 15680
rect 36353 15675 36419 15678
rect 37200 15648 37800 15678
rect 18137 15602 18203 15605
rect 18965 15602 19031 15605
rect 18137 15600 19031 15602
rect 18137 15544 18142 15600
rect 18198 15544 18970 15600
rect 19026 15544 19031 15600
rect 18137 15542 19031 15544
rect 18137 15539 18203 15542
rect 18965 15539 19031 15542
rect 12157 15466 12223 15469
rect 22185 15466 22251 15469
rect 12157 15464 22251 15466
rect 12157 15408 12162 15464
rect 12218 15408 22190 15464
rect 22246 15408 22251 15464
rect 12157 15406 22251 15408
rect 12157 15403 12223 15406
rect 22185 15403 22251 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 200 15058 800 15088
rect 4061 15058 4127 15061
rect 200 15056 4127 15058
rect 200 15000 4066 15056
rect 4122 15000 4127 15056
rect 200 14998 4127 15000
rect 200 14968 800 14998
rect 4061 14995 4127 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 9489 14376 9555 14381
rect 9489 14320 9494 14376
rect 9550 14320 9555 14376
rect 9489 14315 9555 14320
rect 36261 14378 36327 14381
rect 37200 14378 37800 14408
rect 36261 14376 37800 14378
rect 36261 14320 36266 14376
rect 36322 14320 37800 14376
rect 36261 14318 37800 14320
rect 36261 14315 36327 14318
rect 9492 14109 9552 14315
rect 37200 14288 37800 14318
rect 10133 14242 10199 14245
rect 13629 14242 13695 14245
rect 10133 14240 13695 14242
rect 10133 14184 10138 14240
rect 10194 14184 13634 14240
rect 13690 14184 13695 14240
rect 10133 14182 13695 14184
rect 10133 14179 10199 14182
rect 13629 14179 13695 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 9489 14104 9555 14109
rect 9489 14048 9494 14104
rect 9550 14048 9555 14104
rect 9489 14043 9555 14048
rect 10777 13970 10843 13973
rect 18413 13970 18479 13973
rect 10777 13968 18479 13970
rect 10777 13912 10782 13968
rect 10838 13912 18418 13968
rect 18474 13912 18479 13968
rect 10777 13910 18479 13912
rect 10777 13907 10843 13910
rect 18413 13907 18479 13910
rect 10593 13836 10659 13837
rect 10542 13772 10548 13836
rect 10612 13834 10659 13836
rect 10869 13834 10935 13837
rect 10612 13832 10935 13834
rect 10654 13776 10874 13832
rect 10930 13776 10935 13832
rect 10612 13774 10935 13776
rect 10612 13772 10659 13774
rect 10593 13771 10659 13772
rect 10869 13771 10935 13774
rect 200 13698 800 13728
rect 2773 13698 2839 13701
rect 200 13696 2839 13698
rect 200 13640 2778 13696
rect 2834 13640 2839 13696
rect 200 13638 2839 13640
rect 200 13608 800 13638
rect 2773 13635 2839 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 6453 13426 6519 13429
rect 6913 13426 6979 13429
rect 6453 13424 6979 13426
rect 6453 13368 6458 13424
rect 6514 13368 6918 13424
rect 6974 13368 6979 13424
rect 6453 13366 6979 13368
rect 6453 13363 6519 13366
rect 6913 13363 6979 13366
rect 2865 13290 2931 13293
rect 7465 13290 7531 13293
rect 2865 13288 7531 13290
rect 2865 13232 2870 13288
rect 2926 13232 7470 13288
rect 7526 13232 7531 13288
rect 2865 13230 7531 13232
rect 2865 13227 2931 13230
rect 7465 13227 7531 13230
rect 6637 13154 6703 13157
rect 7097 13154 7163 13157
rect 6637 13152 7163 13154
rect 6637 13096 6642 13152
rect 6698 13096 7102 13152
rect 7158 13096 7163 13152
rect 6637 13094 7163 13096
rect 6637 13091 6703 13094
rect 7097 13091 7163 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 3325 13018 3391 13021
rect 8109 13018 8175 13021
rect 3325 13016 8175 13018
rect 3325 12960 3330 13016
rect 3386 12960 8114 13016
rect 8170 12960 8175 13016
rect 3325 12958 8175 12960
rect 3325 12955 3391 12958
rect 8109 12955 8175 12958
rect 6729 12748 6795 12749
rect 6678 12684 6684 12748
rect 6748 12746 6795 12748
rect 6748 12744 6840 12746
rect 6790 12688 6840 12744
rect 6748 12686 6840 12688
rect 6748 12684 6795 12686
rect 6729 12683 6795 12684
rect 6545 12610 6611 12613
rect 8661 12610 8727 12613
rect 6545 12608 8727 12610
rect 6545 12552 6550 12608
rect 6606 12552 8666 12608
rect 8722 12552 8727 12608
rect 6545 12550 8727 12552
rect 6545 12547 6611 12550
rect 8661 12547 8727 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 8477 12474 8543 12477
rect 8937 12474 9003 12477
rect 8477 12472 9003 12474
rect 8477 12416 8482 12472
rect 8538 12416 8942 12472
rect 8998 12416 9003 12472
rect 8477 12414 9003 12416
rect 8477 12411 8543 12414
rect 8937 12411 9003 12414
rect 5349 12338 5415 12341
rect 6545 12338 6611 12341
rect 8661 12338 8727 12341
rect 5349 12336 8727 12338
rect 5349 12280 5354 12336
rect 5410 12280 6550 12336
rect 6606 12280 8666 12336
rect 8722 12280 8727 12336
rect 5349 12278 8727 12280
rect 5349 12275 5415 12278
rect 6545 12275 6611 12278
rect 8661 12275 8727 12278
rect 9857 12338 9923 12341
rect 16113 12338 16179 12341
rect 9857 12336 16179 12338
rect 9857 12280 9862 12336
rect 9918 12280 16118 12336
rect 16174 12280 16179 12336
rect 9857 12278 16179 12280
rect 9857 12275 9923 12278
rect 16113 12275 16179 12278
rect 35801 12338 35867 12341
rect 37200 12338 37800 12368
rect 35801 12336 37800 12338
rect 35801 12280 35806 12336
rect 35862 12280 37800 12336
rect 35801 12278 37800 12280
rect 35801 12275 35867 12278
rect 37200 12248 37800 12278
rect 8109 12202 8175 12205
rect 14457 12202 14523 12205
rect 14917 12202 14983 12205
rect 17217 12202 17283 12205
rect 8109 12200 17283 12202
rect 8109 12144 8114 12200
rect 8170 12144 14462 12200
rect 14518 12144 14922 12200
rect 14978 12144 17222 12200
rect 17278 12144 17283 12200
rect 8109 12142 17283 12144
rect 8109 12139 8175 12142
rect 14457 12139 14523 12142
rect 14917 12139 14983 12142
rect 17217 12139 17283 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 7557 11930 7623 11933
rect 8293 11930 8359 11933
rect 7557 11928 8359 11930
rect 7557 11872 7562 11928
rect 7618 11872 8298 11928
rect 8354 11872 8359 11928
rect 7557 11870 8359 11872
rect 7557 11867 7623 11870
rect 8293 11867 8359 11870
rect 2681 11794 2747 11797
rect 10041 11794 10107 11797
rect 2681 11792 10107 11794
rect 2681 11736 2686 11792
rect 2742 11736 10046 11792
rect 10102 11736 10107 11792
rect 2681 11734 10107 11736
rect 2681 11731 2747 11734
rect 10041 11731 10107 11734
rect 14590 11732 14596 11796
rect 14660 11794 14666 11796
rect 15469 11794 15535 11797
rect 14660 11792 15535 11794
rect 14660 11736 15474 11792
rect 15530 11736 15535 11792
rect 14660 11734 15535 11736
rect 14660 11732 14666 11734
rect 15469 11731 15535 11734
rect 200 11658 800 11688
rect 3785 11658 3851 11661
rect 200 11656 3851 11658
rect 200 11600 3790 11656
rect 3846 11600 3851 11656
rect 200 11598 3851 11600
rect 200 11568 800 11598
rect 3785 11595 3851 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 12709 11386 12775 11389
rect 17401 11386 17467 11389
rect 12709 11384 17467 11386
rect 12709 11328 12714 11384
rect 12770 11328 17406 11384
rect 17462 11328 17467 11384
rect 12709 11326 17467 11328
rect 12709 11323 12775 11326
rect 17401 11323 17467 11326
rect 6361 11250 6427 11253
rect 9489 11250 9555 11253
rect 6361 11248 9555 11250
rect 6361 11192 6366 11248
rect 6422 11192 9494 11248
rect 9550 11192 9555 11248
rect 6361 11190 9555 11192
rect 6361 11187 6427 11190
rect 9489 11187 9555 11190
rect 36261 10978 36327 10981
rect 37200 10978 37800 11008
rect 36261 10976 37800 10978
rect 36261 10920 36266 10976
rect 36322 10920 37800 10976
rect 36261 10918 37800 10920
rect 36261 10915 36327 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 37200 10888 37800 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 3969 10298 4035 10301
rect 200 10296 4035 10298
rect 200 10240 3974 10296
rect 4030 10240 4035 10296
rect 200 10238 4035 10240
rect 200 10208 800 10238
rect 3969 10235 4035 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 7281 9754 7347 9757
rect 8385 9754 8451 9757
rect 7281 9752 8451 9754
rect 7281 9696 7286 9752
rect 7342 9696 8390 9752
rect 8446 9696 8451 9752
rect 7281 9694 8451 9696
rect 7281 9691 7347 9694
rect 8385 9691 8451 9694
rect 1577 9618 1643 9621
rect 4654 9618 4660 9620
rect 1577 9616 4660 9618
rect 1577 9560 1582 9616
rect 1638 9560 4660 9616
rect 1577 9558 4660 9560
rect 1577 9555 1643 9558
rect 4654 9556 4660 9558
rect 4724 9556 4730 9620
rect 7189 9346 7255 9349
rect 9489 9346 9555 9349
rect 7189 9344 9555 9346
rect 7189 9288 7194 9344
rect 7250 9288 9494 9344
rect 9550 9288 9555 9344
rect 7189 9286 9555 9288
rect 7189 9283 7255 9286
rect 9489 9283 9555 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 7465 9210 7531 9213
rect 13997 9210 14063 9213
rect 7465 9208 14063 9210
rect 7465 9152 7470 9208
rect 7526 9152 14002 9208
rect 14058 9152 14063 9208
rect 7465 9150 14063 9152
rect 7465 9147 7531 9150
rect 13997 9147 14063 9150
rect 7925 9074 7991 9077
rect 10726 9074 10732 9076
rect 7925 9072 10732 9074
rect 7925 9016 7930 9072
rect 7986 9016 10732 9072
rect 7925 9014 10732 9016
rect 7925 9011 7991 9014
rect 10726 9012 10732 9014
rect 10796 9012 10802 9076
rect 6085 8938 6151 8941
rect 12341 8938 12407 8941
rect 6085 8936 12407 8938
rect 6085 8880 6090 8936
rect 6146 8880 12346 8936
rect 12402 8880 12407 8936
rect 6085 8878 12407 8880
rect 6085 8875 6151 8878
rect 12341 8875 12407 8878
rect 36261 8938 36327 8941
rect 37200 8938 37800 8968
rect 36261 8936 37800 8938
rect 36261 8880 36266 8936
rect 36322 8880 37800 8936
rect 36261 8878 37800 8880
rect 36261 8875 36327 8878
rect 37200 8848 37800 8878
rect 1945 8802 2011 8805
rect 7373 8802 7439 8805
rect 1945 8800 7439 8802
rect 1945 8744 1950 8800
rect 2006 8744 7378 8800
rect 7434 8744 7439 8800
rect 1945 8742 7439 8744
rect 1945 8739 2011 8742
rect 7373 8739 7439 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 7465 8666 7531 8669
rect 8385 8666 8451 8669
rect 7465 8664 8451 8666
rect 7465 8608 7470 8664
rect 7526 8608 8390 8664
rect 8446 8608 8451 8664
rect 7465 8606 8451 8608
rect 7465 8603 7531 8606
rect 8385 8603 8451 8606
rect 2814 8468 2820 8532
rect 2884 8530 2890 8532
rect 4889 8530 4955 8533
rect 7097 8530 7163 8533
rect 2884 8528 4955 8530
rect 2884 8472 4894 8528
rect 4950 8472 4955 8528
rect 2884 8470 4955 8472
rect 2884 8468 2890 8470
rect 4889 8467 4955 8470
rect 7054 8528 7163 8530
rect 7054 8472 7102 8528
rect 7158 8472 7163 8528
rect 7054 8467 7163 8472
rect 200 8258 800 8288
rect 7054 8261 7114 8467
rect 7649 8394 7715 8397
rect 12433 8394 12499 8397
rect 7649 8392 12499 8394
rect 7649 8336 7654 8392
rect 7710 8336 12438 8392
rect 12494 8336 12499 8392
rect 7649 8334 12499 8336
rect 7649 8331 7715 8334
rect 12433 8331 12499 8334
rect 3969 8258 4035 8261
rect 200 8256 4035 8258
rect 200 8200 3974 8256
rect 4030 8200 4035 8256
rect 200 8198 4035 8200
rect 7054 8256 7163 8261
rect 7054 8200 7102 8256
rect 7158 8200 7163 8256
rect 7054 8198 7163 8200
rect 200 8168 800 8198
rect 3969 8195 4035 8198
rect 7097 8195 7163 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 36261 7578 36327 7581
rect 37200 7578 37800 7608
rect 36261 7576 37800 7578
rect 36261 7520 36266 7576
rect 36322 7520 37800 7576
rect 36261 7518 37800 7520
rect 36261 7515 36327 7518
rect 37200 7488 37800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 2773 6898 2839 6901
rect 200 6896 2839 6898
rect 200 6840 2778 6896
rect 2834 6840 2839 6896
rect 200 6838 2839 6840
rect 200 6808 800 6838
rect 2773 6835 2839 6838
rect 6678 6836 6684 6900
rect 6748 6898 6754 6900
rect 7465 6898 7531 6901
rect 6748 6896 7531 6898
rect 6748 6840 7470 6896
rect 7526 6840 7531 6896
rect 6748 6838 7531 6840
rect 6748 6836 6754 6838
rect 7465 6835 7531 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 2313 5674 2379 5677
rect 10542 5674 10548 5676
rect 2313 5672 10548 5674
rect 2313 5616 2318 5672
rect 2374 5616 10548 5672
rect 2313 5614 10548 5616
rect 2313 5611 2379 5614
rect 10542 5612 10548 5614
rect 10612 5612 10618 5676
rect 15326 5612 15332 5676
rect 15396 5674 15402 5676
rect 35525 5674 35591 5677
rect 15396 5672 35591 5674
rect 15396 5616 35530 5672
rect 35586 5616 35591 5672
rect 15396 5614 35591 5616
rect 15396 5612 15402 5614
rect 35525 5611 35591 5614
rect 36261 5538 36327 5541
rect 37200 5538 37800 5568
rect 36261 5536 37800 5538
rect 36261 5480 36266 5536
rect 36322 5480 37800 5536
rect 36261 5478 37800 5480
rect 36261 5475 36327 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 37200 5448 37800 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1669 4858 1735 4861
rect 200 4856 1735 4858
rect 200 4800 1674 4856
rect 1730 4800 1735 4856
rect 200 4798 1735 4800
rect 200 4768 800 4798
rect 1669 4795 1735 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 36261 4178 36327 4181
rect 37200 4178 37800 4208
rect 36261 4176 37800 4178
rect 36261 4120 36266 4176
rect 36322 4120 37800 4176
rect 36261 4118 37800 4120
rect 36261 4115 36327 4118
rect 37200 4088 37800 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 35801 2138 35867 2141
rect 37200 2138 37800 2168
rect 35801 2136 37800 2138
rect 35801 2080 35806 2136
rect 35862 2080 37800 2136
rect 35801 2078 37800 2080
rect 35801 2075 35867 2078
rect 37200 2048 37800 2078
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 36353 1458 36419 1461
rect 36353 1456 37290 1458
rect 36353 1400 36358 1456
rect 36414 1400 37290 1456
rect 36353 1398 37290 1400
rect 36353 1395 36419 1398
rect 37230 1050 37290 1398
rect 37046 990 37290 1050
rect 37046 778 37106 990
rect 37200 778 37800 808
rect 37046 718 37800 778
rect 37200 688 37800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 1900 36272 1964 36276
rect 1900 36216 1914 36272
rect 1914 36216 1964 36272
rect 1900 36212 1964 36216
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 12572 29472 12636 29476
rect 12572 29416 12586 29472
rect 12586 29416 12636 29472
rect 12572 29412 12636 29416
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 2084 27372 2148 27436
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 12204 25740 12268 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 14596 25060 14660 25124
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 15332 24984 15396 24988
rect 15332 24928 15346 24984
rect 15346 24928 15396 24984
rect 15332 24924 15396 24928
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 2820 23488 2884 23492
rect 2820 23432 2834 23488
rect 2834 23432 2884 23488
rect 2820 23428 2884 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 1900 23156 1964 23220
rect 10732 23080 10796 23084
rect 10732 23024 10746 23080
rect 10746 23024 10796 23080
rect 10732 23020 10796 23024
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 9812 22808 9876 22812
rect 9812 22752 9862 22808
rect 9862 22752 9876 22808
rect 9812 22748 9876 22752
rect 8340 22672 8404 22676
rect 8340 22616 8390 22672
rect 8390 22616 8404 22672
rect 8340 22612 8404 22616
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4660 22068 4724 22132
rect 7972 21796 8036 21860
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 9812 21524 9876 21588
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 12572 20980 12636 21044
rect 8708 20904 8772 20908
rect 8708 20848 8722 20904
rect 8722 20848 8772 20904
rect 8708 20844 8772 20848
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 8340 20572 8404 20636
rect 2084 20300 2148 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 8708 19892 8772 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 7972 19408 8036 19412
rect 7972 19352 8022 19408
rect 8022 19352 8036 19408
rect 7972 19348 8036 19352
rect 4660 19212 4724 19276
rect 12204 19212 12268 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 10548 13832 10612 13836
rect 10548 13776 10598 13832
rect 10598 13776 10612 13832
rect 10548 13772 10612 13776
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 6684 12744 6748 12748
rect 6684 12688 6734 12744
rect 6734 12688 6748 12744
rect 6684 12684 6748 12688
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 14596 11732 14660 11796
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4660 9556 4724 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 10732 9012 10796 9076
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 2820 8468 2884 8532
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 6684 6836 6748 6900
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 10548 5612 10612 5676
rect 15332 5612 15396 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 1899 36276 1965 36277
rect 1899 36212 1900 36276
rect 1964 36212 1965 36276
rect 1899 36211 1965 36212
rect 1902 23221 1962 36211
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 12571 29476 12637 29477
rect 12571 29412 12572 29476
rect 12636 29412 12637 29476
rect 12571 29411 12637 29412
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 2083 27436 2149 27437
rect 2083 27372 2084 27436
rect 2148 27372 2149 27436
rect 2083 27371 2149 27372
rect 1899 23220 1965 23221
rect 1899 23156 1900 23220
rect 1964 23156 1965 23220
rect 1899 23155 1965 23156
rect 2086 20365 2146 27371
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 12203 25804 12269 25805
rect 12203 25740 12204 25804
rect 12268 25740 12269 25804
rect 12203 25739 12269 25740
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 2819 23492 2885 23493
rect 2819 23428 2820 23492
rect 2884 23428 2885 23492
rect 2819 23427 2885 23428
rect 2083 20364 2149 20365
rect 2083 20300 2084 20364
rect 2148 20300 2149 20364
rect 2083 20299 2149 20300
rect 2822 8533 2882 23427
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 10731 23084 10797 23085
rect 10731 23020 10732 23084
rect 10796 23020 10797 23084
rect 10731 23019 10797 23020
rect 9811 22812 9877 22813
rect 9811 22748 9812 22812
rect 9876 22748 9877 22812
rect 9811 22747 9877 22748
rect 8339 22676 8405 22677
rect 8339 22612 8340 22676
rect 8404 22612 8405 22676
rect 8339 22611 8405 22612
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4659 22132 4725 22133
rect 4659 22068 4660 22132
rect 4724 22068 4725 22132
rect 4659 22067 4725 22068
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4662 19277 4722 22067
rect 7971 21860 8037 21861
rect 7971 21796 7972 21860
rect 8036 21796 8037 21860
rect 7971 21795 8037 21796
rect 7974 19413 8034 21795
rect 8342 20637 8402 22611
rect 9814 21589 9874 22747
rect 9811 21588 9877 21589
rect 9811 21524 9812 21588
rect 9876 21524 9877 21588
rect 9811 21523 9877 21524
rect 8707 20908 8773 20909
rect 8707 20844 8708 20908
rect 8772 20844 8773 20908
rect 8707 20843 8773 20844
rect 8339 20636 8405 20637
rect 8339 20572 8340 20636
rect 8404 20572 8405 20636
rect 8339 20571 8405 20572
rect 8710 19957 8770 20843
rect 8707 19956 8773 19957
rect 8707 19892 8708 19956
rect 8772 19892 8773 19956
rect 8707 19891 8773 19892
rect 7971 19412 8037 19413
rect 7971 19348 7972 19412
rect 8036 19348 8037 19412
rect 7971 19347 8037 19348
rect 4659 19276 4725 19277
rect 4659 19212 4660 19276
rect 4724 19212 4725 19276
rect 4659 19211 4725 19212
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4662 9621 4722 19211
rect 10547 13836 10613 13837
rect 10547 13772 10548 13836
rect 10612 13772 10613 13836
rect 10547 13771 10613 13772
rect 6683 12748 6749 12749
rect 6683 12684 6684 12748
rect 6748 12684 6749 12748
rect 6683 12683 6749 12684
rect 4659 9620 4725 9621
rect 4659 9556 4660 9620
rect 4724 9556 4725 9620
rect 4659 9555 4725 9556
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 2819 8532 2885 8533
rect 2819 8468 2820 8532
rect 2884 8468 2885 8532
rect 2819 8467 2885 8468
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 6686 6901 6746 12683
rect 6683 6900 6749 6901
rect 6683 6836 6684 6900
rect 6748 6836 6749 6900
rect 6683 6835 6749 6836
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 10550 5677 10610 13771
rect 10734 9077 10794 23019
rect 12206 19277 12266 25739
rect 12574 21045 12634 29411
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 14595 25124 14661 25125
rect 14595 25060 14596 25124
rect 14660 25060 14661 25124
rect 14595 25059 14661 25060
rect 12571 21044 12637 21045
rect 12571 20980 12572 21044
rect 12636 20980 12637 21044
rect 12571 20979 12637 20980
rect 12203 19276 12269 19277
rect 12203 19212 12204 19276
rect 12268 19212 12269 19276
rect 12203 19211 12269 19212
rect 14598 11797 14658 25059
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 15331 24988 15397 24989
rect 15331 24924 15332 24988
rect 15396 24924 15397 24988
rect 15331 24923 15397 24924
rect 14595 11796 14661 11797
rect 14595 11732 14596 11796
rect 14660 11732 14661 11796
rect 14595 11731 14661 11732
rect 10731 9076 10797 9077
rect 10731 9012 10732 9076
rect 10796 9012 10797 9076
rect 10731 9011 10797 9012
rect 15334 5677 15394 24923
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 10547 5676 10613 5677
rect 10547 5612 10548 5676
rect 10612 5612 10613 5676
rect 10547 5611 10613 5612
rect 15331 5676 15397 5677
rect 15331 5612 15332 5676
rect 15396 5612 15397 5676
rect 15331 5611 15397 5612
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5888 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1667941163
transform -1 0 5244 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1667941163
transform 1 0 4784 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1667941163
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1667941163
transform 1 0 10856 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1667941163
transform -1 0 4140 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1667941163
transform 1 0 10580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1667941163
transform 1 0 11040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1667941163
transform -1 0 9660 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1667941163
transform 1 0 5336 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1667941163
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1667941163
transform 1 0 23000 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1667941163
transform -1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1667941163
transform -1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A
timestamp 1667941163
transform 1 0 20792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1667941163
transform -1 0 24012 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A
timestamp 1667941163
transform -1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1667941163
transform -1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1667941163
transform -1 0 6900 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1667941163
transform 1 0 14536 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1667941163
transform 1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A
timestamp 1667941163
transform 1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1667941163
transform 1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1667941163
transform -1 0 21804 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1667941163
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1667941163
transform 1 0 12696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1667941163
transform -1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform -1 0 18216 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1667941163
transform 1 0 13340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A
timestamp 1667941163
transform 1 0 17296 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1667941163
transform -1 0 18768 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A
timestamp 1667941163
transform -1 0 17664 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1667941163
transform 1 0 18676 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1667941163
transform -1 0 20148 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1667941163
transform 1 0 19044 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1667941163
transform -1 0 15640 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1667941163
transform 1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1667941163
transform 1 0 18032 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1667941163
transform -1 0 20516 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1667941163
transform -1 0 22172 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1667941163
transform -1 0 21620 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1667941163
transform -1 0 23092 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1667941163
transform 1 0 7820 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1667941163
transform -1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A
timestamp 1667941163
transform 1 0 21344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1667941163
transform -1 0 15916 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1667941163
transform 1 0 20976 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1667941163
transform -1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1667941163
transform 1 0 17572 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1667941163
transform 1 0 13616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1667941163
transform -1 0 10580 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1667941163
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A
timestamp 1667941163
transform -1 0 22172 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1667941163
transform -1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1667941163
transform -1 0 21252 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1667941163
transform 1 0 18032 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1667941163
transform -1 0 18308 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform -1 0 19596 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1667941163
transform 1 0 18768 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1667941163
transform 1 0 19688 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform -1 0 12052 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform 1 0 10764 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1667941163
transform -1 0 22724 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1667941163
transform 1 0 9752 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform 1 0 5888 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1667941163
transform 1 0 15456 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1667941163
transform 1 0 6716 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1667941163
transform -1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1667941163
transform -1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1667941163
transform -1 0 15364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1667941163
transform -1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1667941163
transform 1 0 12880 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1667941163
transform 1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1667941163
transform -1 0 21068 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1667941163
transform 1 0 2760 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1667941163
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1667941163
transform -1 0 29440 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1667941163
transform 1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1667941163
transform 1 0 7820 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1667941163
transform 1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1667941163
transform 1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1667941163
transform 1 0 18584 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1667941163
transform 1 0 20148 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1667941163
transform 1 0 9200 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1667941163
transform -1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1667941163
transform -1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1667941163
transform 1 0 16836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1667941163
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1667941163
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1667941163
transform 1 0 28336 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1667941163
transform -1 0 18860 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1667941163
transform 1 0 22632 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1667941163
transform -1 0 17664 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1667941163
transform 1 0 22632 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A
timestamp 1667941163
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__A
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A
timestamp 1667941163
transform 1 0 18032 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__A
timestamp 1667941163
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A
timestamp 1667941163
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__A
timestamp 1667941163
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1667941163
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__A
timestamp 1667941163
transform 1 0 22448 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1667941163
transform -1 0 16284 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A
timestamp 1667941163
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__A
timestamp 1667941163
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__A
timestamp 1667941163
transform 1 0 4140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__A
timestamp 1667941163
transform -1 0 23184 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1667941163
transform -1 0 5428 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1667941163
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__A
timestamp 1667941163
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__A
timestamp 1667941163
transform -1 0 3220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A
timestamp 1667941163
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__A
timestamp 1667941163
transform 1 0 7268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__A
timestamp 1667941163
transform 1 0 10028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__D
timestamp 1667941163
transform -1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__D
timestamp 1667941163
transform -1 0 22908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__D
timestamp 1667941163
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__D
timestamp 1667941163
transform -1 0 6256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__D
timestamp 1667941163
transform -1 0 4784 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__D
timestamp 1667941163
transform -1 0 2944 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__D
timestamp 1667941163
transform -1 0 4784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__D
timestamp 1667941163
transform -1 0 2944 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__536__D
timestamp 1667941163
transform -1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__D
timestamp 1667941163
transform -1 0 7268 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__538__D
timestamp 1667941163
transform -1 0 7912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__D
timestamp 1667941163
transform -1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__D
timestamp 1667941163
transform -1 0 5244 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__D
timestamp 1667941163
transform 1 0 4508 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__D
timestamp 1667941163
transform -1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__D
timestamp 1667941163
transform -1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__D
timestamp 1667941163
transform -1 0 4692 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__D
timestamp 1667941163
transform -1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__D
timestamp 1667941163
transform -1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__D
timestamp 1667941163
transform -1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__D
timestamp 1667941163
transform -1 0 5796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__D
timestamp 1667941163
transform -1 0 7544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__D
timestamp 1667941163
transform -1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__D
timestamp 1667941163
transform -1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__D
timestamp 1667941163
transform -1 0 4692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__595__A
timestamp 1667941163
transform 1 0 35236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__596__A
timestamp 1667941163
transform -1 0 15272 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__A
timestamp 1667941163
transform -1 0 19596 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__A
timestamp 1667941163
transform -1 0 14444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__A
timestamp 1667941163
transform -1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__A
timestamp 1667941163
transform -1 0 20792 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__A
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__A
timestamp 1667941163
transform -1 0 22908 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__A
timestamp 1667941163
transform -1 0 27324 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__608__A
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__A
timestamp 1667941163
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A
timestamp 1667941163
transform 1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__A
timestamp 1667941163
transform 1 0 14812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__615__A
timestamp 1667941163
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__A
timestamp 1667941163
transform -1 0 19596 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__A
timestamp 1667941163
transform -1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__A
timestamp 1667941163
transform -1 0 19688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A
timestamp 1667941163
transform 1 0 12512 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__A
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__A
timestamp 1667941163
transform 1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A
timestamp 1667941163
transform 1 0 21896 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__A
timestamp 1667941163
transform -1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__A
timestamp 1667941163
transform -1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__A
timestamp 1667941163
transform 1 0 27784 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__A
timestamp 1667941163
transform 1 0 8740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__A
timestamp 1667941163
transform -1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__A
timestamp 1667941163
transform 1 0 13800 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__666__A
timestamp 1667941163
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__674__A
timestamp 1667941163
transform -1 0 19320 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__A
timestamp 1667941163
transform 1 0 4508 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__681__A
timestamp 1667941163
transform -1 0 3128 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__688__A
timestamp 1667941163
transform 1 0 3956 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A
timestamp 1667941163
transform -1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__712__A
timestamp 1667941163
transform -1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__746__A
timestamp 1667941163
transform -1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1667941163
transform -1 0 4140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_prog_clk_A
timestamp 1667941163
transform -1 0 5336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_prog_clk_A
timestamp 1667941163
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_prog_clk_A
timestamp 1667941163
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_prog_clk_A
timestamp 1667941163
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_prog_clk_A
timestamp 1667941163
transform -1 0 22632 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_prog_clk_A
timestamp 1667941163
transform 1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_prog_clk_A
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_prog_clk_A
timestamp 1667941163
transform -1 0 4876 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform 1 0 36248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 32568 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 35696 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 35696 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 1748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 15088 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 35696 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 34960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 2392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 2392 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 36432 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 35696 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform 1 0 26496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 35696 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 30452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform 1 0 34224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 2484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 27324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 34960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 35788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 35696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 1748 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 35696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 6808 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 35696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 1748 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 36432 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1667941163
transform -1 0 35696 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output46_A
timestamp 1667941163
transform 1 0 35512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp 1667941163
transform 1 0 3128 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output50_A
timestamp 1667941163
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1667941163
transform -1 0 22908 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output58_A
timestamp 1667941163
transform 1 0 34960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1667941163
transform 1 0 13800 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1667941163
transform -1 0 2116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1667941163
transform 1 0 35512 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1667941163
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77
timestamp 1667941163
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1667941163
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10120 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1667941163
transform 1 0 10856 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127
timestamp 1667941163
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132
timestamp 1667941163
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_152
timestamp 1667941163
transform 1 0 15088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1667941163
transform 1 0 15824 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1667941163
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_182 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_203
timestamp 1667941163
transform 1 0 19780 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_211
timestamp 1667941163
transform 1 0 20516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1667941163
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1667941163
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_259
timestamp 1667941163
transform 1 0 24932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_267
timestamp 1667941163
transform 1 0 25668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1667941163
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_303
timestamp 1667941163
transform 1 0 28980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_323
timestamp 1667941163
transform 1 0 30820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_331
timestamp 1667941163
transform 1 0 31556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1667941163
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_378
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_384
timestamp 1667941163
transform 1 0 36432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1667941163
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1667941163
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_70
timestamp 1667941163
transform 1 0 7544 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_82
timestamp 1667941163
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 1667941163
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1667941163
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1667941163
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_285
timestamp 1667941163
transform 1 0 27324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_297
timestamp 1667941163
transform 1 0 28428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_309
timestamp 1667941163
transform 1 0 29532 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_319
timestamp 1667941163
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1667941163
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_365
timestamp 1667941163
transform 1 0 34684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1667941163
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_376
timestamp 1667941163
transform 1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_384
timestamp 1667941163
transform 1 0 36432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_214
timestamp 1667941163
transform 1 0 20792 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_226
timestamp 1667941163
transform 1 0 21896 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_238
timestamp 1667941163
transform 1 0 23000 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_373
timestamp 1667941163
transform 1 0 35420 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_376
timestamp 1667941163
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_384
timestamp 1667941163
transform 1 0 36432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_10
timestamp 1667941163
transform 1 0 2024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_17
timestamp 1667941163
transform 1 0 2668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_23
timestamp 1667941163
transform 1 0 3220 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_31
timestamp 1667941163
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_43
timestamp 1667941163
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1667941163
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_12
timestamp 1667941163
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_23
timestamp 1667941163
transform 1 0 3220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_33
timestamp 1667941163
transform 1 0 4140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp 1667941163
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_40
timestamp 1667941163
transform 1 0 4784 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_46
timestamp 1667941163
transform 1 0 5336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_58
timestamp 1667941163
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1667941163
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_90
timestamp 1667941163
transform 1 0 9384 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_102
timestamp 1667941163
transform 1 0 10488 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_114
timestamp 1667941163
transform 1 0 11592 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_126
timestamp 1667941163
transform 1 0 12696 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_384
timestamp 1667941163
transform 1 0 36432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_19
timestamp 1667941163
transform 1 0 2852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_26
timestamp 1667941163
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_175
timestamp 1667941163
transform 1 0 17204 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1667941163
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1667941163
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1667941163
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1667941163
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_46
timestamp 1667941163
transform 1 0 5336 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_56
timestamp 1667941163
transform 1 0 6256 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1667941163
transform 1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_66
timestamp 1667941163
transform 1 0 7176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_69
timestamp 1667941163
transform 1 0 7452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1667941163
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_373
timestamp 1667941163
transform 1 0 35420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_376
timestamp 1667941163
transform 1 0 35696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_384
timestamp 1667941163
transform 1 0 36432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_26
timestamp 1667941163
transform 1 0 3496 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_32
timestamp 1667941163
transform 1 0 4048 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1667941163
transform 1 0 4416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_43
timestamp 1667941163
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_61
timestamp 1667941163
transform 1 0 6716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_67
timestamp 1667941163
transform 1 0 7268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1667941163
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_74
timestamp 1667941163
transform 1 0 7912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_77
timestamp 1667941163
transform 1 0 8188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_87
timestamp 1667941163
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_99
timestamp 1667941163
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_130
timestamp 1667941163
transform 1 0 13064 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_142
timestamp 1667941163
transform 1 0 14168 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_154
timestamp 1667941163
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_231
timestamp 1667941163
transform 1 0 22356 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_33
timestamp 1667941163
transform 1 0 4140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1667941163
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_47
timestamp 1667941163
transform 1 0 5428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_54
timestamp 1667941163
transform 1 0 6072 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_62
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_71
timestamp 1667941163
transform 1 0 7636 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_79
timestamp 1667941163
transform 1 0 8372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_89
timestamp 1667941163
transform 1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1667941163
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1667941163
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_102
timestamp 1667941163
transform 1 0 10488 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_110
timestamp 1667941163
transform 1 0 11224 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_122
timestamp 1667941163
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp 1667941163
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_229
timestamp 1667941163
transform 1 0 22172 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_234
timestamp 1667941163
transform 1 0 22632 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1667941163
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_385
timestamp 1667941163
transform 1 0 36524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_25
timestamp 1667941163
transform 1 0 3404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1667941163
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1667941163
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_68
timestamp 1667941163
transform 1 0 7360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1667941163
transform 1 0 7912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_87
timestamp 1667941163
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_94
timestamp 1667941163
transform 1 0 9752 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1667941163
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_119
timestamp 1667941163
transform 1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_71
timestamp 1667941163
transform 1 0 7636 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1667941163
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_96
timestamp 1667941163
transform 1 0 9936 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1667941163
transform 1 0 10672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1667941163
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1667941163
transform 1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_119
timestamp 1667941163
transform 1 0 12052 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1667941163
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1667941163
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_132
timestamp 1667941163
transform 1 0 13248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1667941163
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_373
timestamp 1667941163
transform 1 0 35420 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_376
timestamp 1667941163
transform 1 0 35696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_384
timestamp 1667941163
transform 1 0 36432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_12
timestamp 1667941163
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_36
timestamp 1667941163
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_43
timestamp 1667941163
transform 1 0 5060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1667941163
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_63
timestamp 1667941163
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1667941163
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1667941163
transform 1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1667941163
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1667941163
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_104
timestamp 1667941163
transform 1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_118
timestamp 1667941163
transform 1 0 11960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_128
timestamp 1667941163
transform 1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_132
timestamp 1667941163
transform 1 0 13248 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_135
timestamp 1667941163
transform 1 0 13524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_139
timestamp 1667941163
transform 1 0 13892 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1667941163
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_148
timestamp 1667941163
transform 1 0 14720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1667941163
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_174
timestamp 1667941163
transform 1 0 17112 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_186
timestamp 1667941163
transform 1 0 18216 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_198
timestamp 1667941163
transform 1 0 19320 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_210
timestamp 1667941163
transform 1 0 20424 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1667941163
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_33
timestamp 1667941163
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_54
timestamp 1667941163
transform 1 0 6072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1667941163
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_68
timestamp 1667941163
transform 1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1667941163
transform 1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1667941163
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_101
timestamp 1667941163
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_108
timestamp 1667941163
transform 1 0 11040 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1667941163
transform 1 0 11776 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1667941163
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1667941163
transform 1 0 12788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_145
timestamp 1667941163
transform 1 0 14444 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_151
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_157
timestamp 1667941163
transform 1 0 15548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_169
timestamp 1667941163
transform 1 0 16652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_181
timestamp 1667941163
transform 1 0 17756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1667941163
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_373
timestamp 1667941163
transform 1 0 35420 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_376
timestamp 1667941163
transform 1 0 35696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_384
timestamp 1667941163
transform 1 0 36432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_25
timestamp 1667941163
transform 1 0 3404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_33
timestamp 1667941163
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_79
timestamp 1667941163
transform 1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1667941163
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_92
timestamp 1667941163
transform 1 0 9568 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_98
timestamp 1667941163
transform 1 0 10120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1667941163
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1667941163
transform 1 0 12420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_130
timestamp 1667941163
transform 1 0 13064 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_136
timestamp 1667941163
transform 1 0 13616 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_140
timestamp 1667941163
transform 1 0 13984 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_151
timestamp 1667941163
transform 1 0 14996 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1667941163
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_35
timestamp 1667941163
transform 1 0 4324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_43
timestamp 1667941163
transform 1 0 5060 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_49
timestamp 1667941163
transform 1 0 5612 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_71
timestamp 1667941163
transform 1 0 7636 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_91
timestamp 1667941163
transform 1 0 9476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_95
timestamp 1667941163
transform 1 0 9844 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1667941163
transform 1 0 10488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_108
timestamp 1667941163
transform 1 0 11040 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1667941163
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_152
timestamp 1667941163
transform 1 0 15088 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp 1667941163
transform 1 0 15640 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1667941163
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_168
timestamp 1667941163
transform 1 0 16560 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_174
timestamp 1667941163
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_186
timestamp 1667941163
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_385
timestamp 1667941163
transform 1 0 36524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1667941163
transform 1 0 2208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1667941163
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_43
timestamp 1667941163
transform 1 0 5060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 1667941163
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1667941163
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_100
timestamp 1667941163
transform 1 0 10304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1667941163
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_124
timestamp 1667941163
transform 1 0 12512 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 1667941163
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_138
timestamp 1667941163
transform 1 0 13800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_151
timestamp 1667941163
transform 1 0 14996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_155
timestamp 1667941163
transform 1 0 15364 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1667941163
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_180
timestamp 1667941163
transform 1 0 17664 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1667941163
transform 1 0 18768 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1667941163
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_202
timestamp 1667941163
transform 1 0 19688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214
timestamp 1667941163
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1667941163
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1667941163
transform 1 0 6072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_58
timestamp 1667941163
transform 1 0 6440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_108
timestamp 1667941163
transform 1 0 11040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_118
timestamp 1667941163
transform 1 0 11960 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_124
timestamp 1667941163
transform 1 0 12512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 1667941163
transform 1 0 12880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1667941163
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 1667941163
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1667941163
transform 1 0 17480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1667941163
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_201
timestamp 1667941163
transform 1 0 19596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_213
timestamp 1667941163
transform 1 0 20700 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_225
timestamp 1667941163
transform 1 0 21804 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_237
timestamp 1667941163
transform 1 0 22908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1667941163
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_384
timestamp 1667941163
transform 1 0 36432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_25
timestamp 1667941163
transform 1 0 3404 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_63
timestamp 1667941163
transform 1 0 6900 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_92
timestamp 1667941163
transform 1 0 9568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_96
timestamp 1667941163
transform 1 0 9936 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_100
timestamp 1667941163
transform 1 0 10304 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_121
timestamp 1667941163
transform 1 0 12236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_128
timestamp 1667941163
transform 1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_135
timestamp 1667941163
transform 1 0 13524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_141
timestamp 1667941163
transform 1 0 14076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1667941163
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1667941163
transform 1 0 15088 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1667941163
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1667941163
transform 1 0 18032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_191
timestamp 1667941163
transform 1 0 18676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1667941163
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1667941163
transform 1 0 19872 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_210
timestamp 1667941163
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1667941163
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_33
timestamp 1667941163
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1667941163
transform 1 0 6072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_58
timestamp 1667941163
transform 1 0 6440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1667941163
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1667941163
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1667941163
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1667941163
transform 1 0 11960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_122
timestamp 1667941163
transform 1 0 12328 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_132
timestamp 1667941163
transform 1 0 13248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_146
timestamp 1667941163
transform 1 0 14536 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_159
timestamp 1667941163
transform 1 0 15732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_167
timestamp 1667941163
transform 1 0 16468 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_171
timestamp 1667941163
transform 1 0 16836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_184
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1667941163
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_216
timestamp 1667941163
transform 1 0 20976 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_228
timestamp 1667941163
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_240
timestamp 1667941163
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_385
timestamp 1667941163
transform 1 0 36524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1667941163
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1667941163
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_63
timestamp 1667941163
transform 1 0 6900 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_90
timestamp 1667941163
transform 1 0 9384 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_94
timestamp 1667941163
transform 1 0 9752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1667941163
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1667941163
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1667941163
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_151
timestamp 1667941163
transform 1 0 14996 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1667941163
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_186
timestamp 1667941163
transform 1 0 18216 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_192
timestamp 1667941163
transform 1 0 18768 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1667941163
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1667941163
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_216
timestamp 1667941163
transform 1 0 20976 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_229
timestamp 1667941163
transform 1 0 22172 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_241
timestamp 1667941163
transform 1 0 23276 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_253
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_265
timestamp 1667941163
transform 1 0 25484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1667941163
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_376
timestamp 1667941163
transform 1 0 35696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_384
timestamp 1667941163
transform 1 0 36432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_55
timestamp 1667941163
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_89
timestamp 1667941163
transform 1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1667941163
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_103
timestamp 1667941163
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_111
timestamp 1667941163
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1667941163
transform 1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_128
timestamp 1667941163
transform 1 0 12880 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_134
timestamp 1667941163
transform 1 0 13432 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1667941163
transform 1 0 14720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_155
timestamp 1667941163
transform 1 0 15364 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1667941163
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_179
timestamp 1667941163
transform 1 0 17572 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1667941163
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1667941163
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_201
timestamp 1667941163
transform 1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_205
timestamp 1667941163
transform 1 0 19964 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1667941163
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_216
timestamp 1667941163
transform 1 0 20976 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1667941163
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_234
timestamp 1667941163
transform 1 0 22632 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1667941163
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_381
timestamp 1667941163
transform 1 0 36156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_385
timestamp 1667941163
transform 1 0 36524 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_26
timestamp 1667941163
transform 1 0 3496 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_61
timestamp 1667941163
transform 1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_88
timestamp 1667941163
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1667941163
transform 1 0 10028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1667941163
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_117
timestamp 1667941163
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_121
timestamp 1667941163
transform 1 0 12236 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_134
timestamp 1667941163
transform 1 0 13432 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_140
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_150
timestamp 1667941163
transform 1 0 14904 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1667941163
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1667941163
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_202
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_212
timestamp 1667941163
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1667941163
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_236
timestamp 1667941163
transform 1 0 22816 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_243
timestamp 1667941163
transform 1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_55
timestamp 1667941163
transform 1 0 6164 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1667941163
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_127
timestamp 1667941163
transform 1 0 12788 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1667941163
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1667941163
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_164
timestamp 1667941163
transform 1 0 16192 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1667941163
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_188
timestamp 1667941163
transform 1 0 18400 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 1667941163
transform 1 0 19780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1667941163
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_226
timestamp 1667941163
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_239
timestamp 1667941163
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_373
timestamp 1667941163
transform 1 0 35420 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_376
timestamp 1667941163
transform 1 0 35696 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_384
timestamp 1667941163
transform 1 0 36432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_28
timestamp 1667941163
transform 1 0 3680 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1667941163
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1667941163
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_66
timestamp 1667941163
transform 1 0 7176 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_90
timestamp 1667941163
transform 1 0 9384 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1667941163
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1667941163
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_118
timestamp 1667941163
transform 1 0 11960 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_126
timestamp 1667941163
transform 1 0 12696 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 1667941163
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1667941163
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1667941163
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1667941163
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_200
timestamp 1667941163
transform 1 0 19504 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1667941163
transform 1 0 20700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1667941163
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_229
timestamp 1667941163
transform 1 0 22172 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_235
timestamp 1667941163
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_247
timestamp 1667941163
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_259
timestamp 1667941163
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1667941163
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1667941163
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 1667941163
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1667941163
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_108
timestamp 1667941163
transform 1 0 11040 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1667941163
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_147
timestamp 1667941163
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_151
timestamp 1667941163
transform 1 0 14996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_164
timestamp 1667941163
transform 1 0 16192 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_171
timestamp 1667941163
transform 1 0 16836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1667941163
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1667941163
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_203
timestamp 1667941163
transform 1 0 19780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1667941163
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_225
timestamp 1667941163
transform 1 0 21804 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_231
timestamp 1667941163
transform 1 0 22356 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_237
timestamp 1667941163
transform 1 0 22908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1667941163
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_385
timestamp 1667941163
transform 1 0 36524 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_42
timestamp 1667941163
transform 1 0 4968 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_50
timestamp 1667941163
transform 1 0 5704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_64
timestamp 1667941163
transform 1 0 6992 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_91
timestamp 1667941163
transform 1 0 9476 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_101
timestamp 1667941163
transform 1 0 10396 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_119
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_126
timestamp 1667941163
transform 1 0 12696 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_139
timestamp 1667941163
transform 1 0 13892 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_156
timestamp 1667941163
transform 1 0 15456 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_160
timestamp 1667941163
transform 1 0 15824 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1667941163
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1667941163
transform 1 0 17112 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1667941163
transform 1 0 17848 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1667941163
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_205
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_211
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1667941163
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_229
timestamp 1667941163
transform 1 0 22172 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_235
timestamp 1667941163
transform 1 0 22724 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_247
timestamp 1667941163
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_259
timestamp 1667941163
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_271
timestamp 1667941163
transform 1 0 26036 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1667941163
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_377
timestamp 1667941163
transform 1 0 35788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_384
timestamp 1667941163
transform 1 0 36432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1667941163
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_35
timestamp 1667941163
transform 1 0 4324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp 1667941163
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1667941163
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1667941163
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1667941163
transform 1 0 10948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1667941163
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 1667941163
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_150
timestamp 1667941163
transform 1 0 14904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_163
timestamp 1667941163
transform 1 0 16100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_169
timestamp 1667941163
transform 1 0 16652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_179
timestamp 1667941163
transform 1 0 17572 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_185
timestamp 1667941163
transform 1 0 18124 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_201
timestamp 1667941163
transform 1 0 19596 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_207
timestamp 1667941163
transform 1 0 20148 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_216
timestamp 1667941163
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1667941163
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1667941163
transform 1 0 22080 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_234
timestamp 1667941163
transform 1 0 22632 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1667941163
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_385
timestamp 1667941163
transform 1 0 36524 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1667941163
transform 1 0 2668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_42
timestamp 1667941163
transform 1 0 4968 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_50
timestamp 1667941163
transform 1 0 5704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_63
timestamp 1667941163
transform 1 0 6900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_90
timestamp 1667941163
transform 1 0 9384 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_98
timestamp 1667941163
transform 1 0 10120 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_102
timestamp 1667941163
transform 1 0 10488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_106
timestamp 1667941163
transform 1 0 10856 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1667941163
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1667941163
transform 1 0 14076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1667941163
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_158
timestamp 1667941163
transform 1 0 15640 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1667941163
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_173
timestamp 1667941163
transform 1 0 17020 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_179
timestamp 1667941163
transform 1 0 17572 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_182
timestamp 1667941163
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_189
timestamp 1667941163
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_197
timestamp 1667941163
transform 1 0 19228 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_201
timestamp 1667941163
transform 1 0 19596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_204
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1667941163
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_229
timestamp 1667941163
transform 1 0 22172 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_241
timestamp 1667941163
transform 1 0 23276 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_253
timestamp 1667941163
transform 1 0 24380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_265
timestamp 1667941163
transform 1 0 25484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1667941163
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1667941163
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_35
timestamp 1667941163
transform 1 0 4324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_57
timestamp 1667941163
transform 1 0 6348 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_89
timestamp 1667941163
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1667941163
transform 1 0 9660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_100
timestamp 1667941163
transform 1 0 10304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_107
timestamp 1667941163
transform 1 0 10948 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_111
timestamp 1667941163
transform 1 0 11316 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1667941163
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_158
timestamp 1667941163
transform 1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1667941163
transform 1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_178
timestamp 1667941163
transform 1 0 17480 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_186
timestamp 1667941163
transform 1 0 18216 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_202
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_210
timestamp 1667941163
transform 1 0 20424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_220
timestamp 1667941163
transform 1 0 21344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_224
timestamp 1667941163
transform 1 0 21712 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1667941163
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_234
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_240
timestamp 1667941163
transform 1 0 23184 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_385
timestamp 1667941163
transform 1 0 36524 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_29
timestamp 1667941163
transform 1 0 3772 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1667941163
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_62
timestamp 1667941163
transform 1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_89
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_97
timestamp 1667941163
transform 1 0 10028 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_101
timestamp 1667941163
transform 1 0 10396 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_126
timestamp 1667941163
transform 1 0 12696 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_134
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1667941163
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_174
timestamp 1667941163
transform 1 0 17112 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_180
timestamp 1667941163
transform 1 0 17664 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_183
timestamp 1667941163
transform 1 0 17940 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_192
timestamp 1667941163
transform 1 0 18768 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1667941163
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_214
timestamp 1667941163
transform 1 0 20792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1667941163
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_229
timestamp 1667941163
transform 1 0 22172 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_233
timestamp 1667941163
transform 1 0 22540 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_239
timestamp 1667941163
transform 1 0 23092 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_251
timestamp 1667941163
transform 1 0 24196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_260
timestamp 1667941163
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_266
timestamp 1667941163
transform 1 0 25576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_379
timestamp 1667941163
transform 1 0 35972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_384
timestamp 1667941163
transform 1 0 36432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_54
timestamp 1667941163
transform 1 0 6072 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1667941163
transform 1 0 9292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1667941163
transform 1 0 9660 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_100
timestamp 1667941163
transform 1 0 10304 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_107
timestamp 1667941163
transform 1 0 10948 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1667941163
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_145
timestamp 1667941163
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_158
timestamp 1667941163
transform 1 0 15640 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_167
timestamp 1667941163
transform 1 0 16468 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1667941163
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1667941163
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_212
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_227
timestamp 1667941163
transform 1 0 21988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_239
timestamp 1667941163
transform 1 0 23092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_385
timestamp 1667941163
transform 1 0 36524 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_28
timestamp 1667941163
transform 1 0 3680 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1667941163
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_65
timestamp 1667941163
transform 1 0 7084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_92
timestamp 1667941163
transform 1 0 9568 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1667941163
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_119
timestamp 1667941163
transform 1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1667941163
transform 1 0 13248 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_138
timestamp 1667941163
transform 1 0 13800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1667941163
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_152
timestamp 1667941163
transform 1 0 15088 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1667941163
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_180
timestamp 1667941163
transform 1 0 17664 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1667941163
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_202
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1667941163
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1667941163
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_236
timestamp 1667941163
transform 1 0 22816 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_248
timestamp 1667941163
transform 1 0 23920 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_260
timestamp 1667941163
transform 1 0 25024 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_272
timestamp 1667941163
transform 1 0 26128 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_377
timestamp 1667941163
transform 1 0 35788 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_381
timestamp 1667941163
transform 1 0 36156 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_33
timestamp 1667941163
transform 1 0 4140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_54
timestamp 1667941163
transform 1 0 6072 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_60
timestamp 1667941163
transform 1 0 6624 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_104
timestamp 1667941163
transform 1 0 10672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_111
timestamp 1667941163
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_124
timestamp 1667941163
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1667941163
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1667941163
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_150
timestamp 1667941163
transform 1 0 14904 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1667941163
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1667941163
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1667941163
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1667941163
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1667941163
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1667941163
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_191
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_208
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_220
timestamp 1667941163
transform 1 0 21344 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_228
timestamp 1667941163
transform 1 0 22080 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_239
timestamp 1667941163
transform 1 0 23092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_385
timestamp 1667941163
transform 1 0 36524 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_26
timestamp 1667941163
transform 1 0 3496 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_63
timestamp 1667941163
transform 1 0 6900 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_90
timestamp 1667941163
transform 1 0 9384 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1667941163
transform 1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1667941163
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_122
timestamp 1667941163
transform 1 0 12328 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1667941163
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_148
timestamp 1667941163
transform 1 0 14720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_155
timestamp 1667941163
transform 1 0 15364 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1667941163
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_173
timestamp 1667941163
transform 1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1667941163
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1667941163
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1667941163
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_198
timestamp 1667941163
transform 1 0 19320 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_206
timestamp 1667941163
transform 1 0 20056 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_210
timestamp 1667941163
transform 1 0 20424 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1667941163
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_369
timestamp 1667941163
transform 1 0 35052 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_380
timestamp 1667941163
transform 1 0 36064 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_55
timestamp 1667941163
transform 1 0 6164 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1667941163
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_95
timestamp 1667941163
transform 1 0 9844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_102
timestamp 1667941163
transform 1 0 10488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_116
timestamp 1667941163
transform 1 0 11776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_123
timestamp 1667941163
transform 1 0 12420 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1667941163
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_147
timestamp 1667941163
transform 1 0 14628 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_160
timestamp 1667941163
transform 1 0 15824 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_167
timestamp 1667941163
transform 1 0 16468 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_174
timestamp 1667941163
transform 1 0 17112 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_180
timestamp 1667941163
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_186
timestamp 1667941163
transform 1 0 18216 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1667941163
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_208
timestamp 1667941163
transform 1 0 20240 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_220
timestamp 1667941163
transform 1 0 21344 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_232
timestamp 1667941163
transform 1 0 22448 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1667941163
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_385
timestamp 1667941163
transform 1 0 36524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_17
timestamp 1667941163
transform 1 0 2668 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_20
timestamp 1667941163
transform 1 0 2944 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_47
timestamp 1667941163
transform 1 0 5428 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_63
timestamp 1667941163
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_90
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1667941163
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_106
timestamp 1667941163
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_120
timestamp 1667941163
transform 1 0 12144 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1667941163
transform 1 0 12788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_140
timestamp 1667941163
transform 1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_153
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_174
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_178
timestamp 1667941163
transform 1 0 17480 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1667941163
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_376
timestamp 1667941163
transform 1 0 35696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_384
timestamp 1667941163
transform 1 0 36432 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_17
timestamp 1667941163
transform 1 0 2668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_20
timestamp 1667941163
transform 1 0 2944 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_51
timestamp 1667941163
transform 1 0 5796 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_55
timestamp 1667941163
transform 1 0 6164 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_76
timestamp 1667941163
transform 1 0 8096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_91
timestamp 1667941163
transform 1 0 9476 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1667941163
transform 1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_105
timestamp 1667941163
transform 1 0 10764 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_112
timestamp 1667941163
transform 1 0 11408 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1667941163
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1667941163
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_152
timestamp 1667941163
transform 1 0 15088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_159
timestamp 1667941163
transform 1 0 15732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_167
timestamp 1667941163
transform 1 0 16468 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_183
timestamp 1667941163
transform 1 0 17940 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1667941163
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_208
timestamp 1667941163
transform 1 0 20240 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_214
timestamp 1667941163
transform 1 0 20792 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_226
timestamp 1667941163
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_238
timestamp 1667941163
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1667941163
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_271
timestamp 1667941163
transform 1 0 26036 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_275
timestamp 1667941163
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1667941163
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_299
timestamp 1667941163
transform 1 0 28612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_385
timestamp 1667941163
transform 1 0 36524 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_42
timestamp 1667941163
transform 1 0 4968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_48
timestamp 1667941163
transform 1 0 5520 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_63
timestamp 1667941163
transform 1 0 6900 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_67
timestamp 1667941163
transform 1 0 7268 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_92
timestamp 1667941163
transform 1 0 9568 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_103
timestamp 1667941163
transform 1 0 10580 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1667941163
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_131
timestamp 1667941163
transform 1 0 13156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_138
timestamp 1667941163
transform 1 0 13800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_142
timestamp 1667941163
transform 1 0 14168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_152
timestamp 1667941163
transform 1 0 15088 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_158
timestamp 1667941163
transform 1 0 15640 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1667941163
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_180
timestamp 1667941163
transform 1 0 17664 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_187
timestamp 1667941163
transform 1 0 18308 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_199
timestamp 1667941163
transform 1 0 19412 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_203
timestamp 1667941163
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_209
timestamp 1667941163
transform 1 0 20332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 1667941163
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_302
timestamp 1667941163
transform 1 0 28888 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_308
timestamp 1667941163
transform 1 0 29440 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_320
timestamp 1667941163
transform 1 0 30544 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1667941163
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_379
timestamp 1667941163
transform 1 0 35972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_384
timestamp 1667941163
transform 1 0 36432 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_9
timestamp 1667941163
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1667941163
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_20
timestamp 1667941163
transform 1 0 2944 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1667941163
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_33
timestamp 1667941163
transform 1 0 4140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_39
timestamp 1667941163
transform 1 0 4692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_45
timestamp 1667941163
transform 1 0 5244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_69
timestamp 1667941163
transform 1 0 7452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_75
timestamp 1667941163
transform 1 0 8004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_89
timestamp 1667941163
transform 1 0 9292 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1667941163
transform 1 0 9660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_100
timestamp 1667941163
transform 1 0 10304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1667941163
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_120
timestamp 1667941163
transform 1 0 12144 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_128
timestamp 1667941163
transform 1 0 12880 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1667941163
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_160
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_166
timestamp 1667941163
transform 1 0 16376 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1667941163
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_184
timestamp 1667941163
transform 1 0 18032 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_208
timestamp 1667941163
transform 1 0 20240 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_220
timestamp 1667941163
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_232
timestamp 1667941163
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1667941163
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_257
timestamp 1667941163
transform 1 0 24748 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_269
timestamp 1667941163
transform 1 0 25852 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_281
timestamp 1667941163
transform 1 0 26956 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_293
timestamp 1667941163
transform 1 0 28060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1667941163
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_385
timestamp 1667941163
transform 1 0 36524 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_9
timestamp 1667941163
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_13
timestamp 1667941163
transform 1 0 2300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_20
timestamp 1667941163
transform 1 0 2944 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1667941163
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_38
timestamp 1667941163
transform 1 0 4600 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_41
timestamp 1667941163
transform 1 0 4876 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_66
timestamp 1667941163
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_79
timestamp 1667941163
transform 1 0 8372 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_92
timestamp 1667941163
transform 1 0 9568 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_100
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1667941163
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_129
timestamp 1667941163
transform 1 0 12972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_136
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_148
timestamp 1667941163
transform 1 0 14720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_156
timestamp 1667941163
transform 1 0 15456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_180
timestamp 1667941163
transform 1 0 17664 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_191
timestamp 1667941163
transform 1 0 18676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_198
timestamp 1667941163
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_211
timestamp 1667941163
transform 1 0 20516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_236
timestamp 1667941163
transform 1 0 22816 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_248
timestamp 1667941163
transform 1 0 23920 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_260
timestamp 1667941163
transform 1 0 25024 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1667941163
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_287
timestamp 1667941163
transform 1 0 27508 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_291
timestamp 1667941163
transform 1 0 27876 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_297
timestamp 1667941163
transform 1 0 28428 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_309
timestamp 1667941163
transform 1 0 29532 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_321
timestamp 1667941163
transform 1 0 30636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1667941163
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_7
timestamp 1667941163
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_14
timestamp 1667941163
transform 1 0 2392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1667941163
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1667941163
transform 1 0 4784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_47
timestamp 1667941163
transform 1 0 5428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_55
timestamp 1667941163
transform 1 0 6164 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_59
timestamp 1667941163
transform 1 0 6532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_66
timestamp 1667941163
transform 1 0 7176 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_75
timestamp 1667941163
transform 1 0 8004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1667941163
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1667941163
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1667941163
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_112
timestamp 1667941163
transform 1 0 11408 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_125
timestamp 1667941163
transform 1 0 12604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1667941163
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1667941163
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_171
timestamp 1667941163
transform 1 0 16836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_178
timestamp 1667941163
transform 1 0 17480 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1667941163
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_203
timestamp 1667941163
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_207
timestamp 1667941163
transform 1 0 20148 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1667941163
transform 1 0 20700 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_217
timestamp 1667941163
transform 1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_223
timestamp 1667941163
transform 1 0 21620 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_235
timestamp 1667941163
transform 1 0 22724 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1667941163
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_381
timestamp 1667941163
transform 1 0 36156 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_384
timestamp 1667941163
transform 1 0 36432 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_14
timestamp 1667941163
transform 1 0 2392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_20
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_33
timestamp 1667941163
transform 1 0 4140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_47
timestamp 1667941163
transform 1 0 5428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1667941163
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_62
timestamp 1667941163
transform 1 0 6808 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_71
timestamp 1667941163
transform 1 0 7636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_78
timestamp 1667941163
transform 1 0 8280 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_85
timestamp 1667941163
transform 1 0 8924 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_92
timestamp 1667941163
transform 1 0 9568 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1667941163
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_130
timestamp 1667941163
transform 1 0 13064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_143
timestamp 1667941163
transform 1 0 14260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_160
timestamp 1667941163
transform 1 0 15824 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_184
timestamp 1667941163
transform 1 0 18032 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_191
timestamp 1667941163
transform 1 0 18676 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_197
timestamp 1667941163
transform 1 0 19228 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_201
timestamp 1667941163
transform 1 0 19596 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_204
timestamp 1667941163
transform 1 0 19872 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1667941163
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_384
timestamp 1667941163
transform 1 0 36432 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_7
timestamp 1667941163
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_17
timestamp 1667941163
transform 1 0 2668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1667941163
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_33
timestamp 1667941163
transform 1 0 4140 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_39
timestamp 1667941163
transform 1 0 4692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_45
timestamp 1667941163
transform 1 0 5244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_58
timestamp 1667941163
transform 1 0 6440 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_71
timestamp 1667941163
transform 1 0 7636 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_79
timestamp 1667941163
transform 1 0 8372 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_90
timestamp 1667941163
transform 1 0 9384 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_103
timestamp 1667941163
transform 1 0 10580 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_113
timestamp 1667941163
transform 1 0 11500 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_127
timestamp 1667941163
transform 1 0 12788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_147
timestamp 1667941163
transform 1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_151
timestamp 1667941163
transform 1 0 14996 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_156
timestamp 1667941163
transform 1 0 15456 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_164
timestamp 1667941163
transform 1 0 16192 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_188
timestamp 1667941163
transform 1 0 18400 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_201
timestamp 1667941163
transform 1 0 19596 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_207
timestamp 1667941163
transform 1 0 20148 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_217
timestamp 1667941163
transform 1 0 21068 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_229
timestamp 1667941163
transform 1 0 22172 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_241
timestamp 1667941163
transform 1 0 23276 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1667941163
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_385
timestamp 1667941163
transform 1 0 36524 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_14
timestamp 1667941163
transform 1 0 2392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_21
timestamp 1667941163
transform 1 0 3036 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_28
timestamp 1667941163
transform 1 0 3680 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_40
timestamp 1667941163
transform 1 0 4784 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1667941163
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_67
timestamp 1667941163
transform 1 0 7268 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_75
timestamp 1667941163
transform 1 0 8004 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_79
timestamp 1667941163
transform 1 0 8372 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_83
timestamp 1667941163
transform 1 0 8740 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_87
timestamp 1667941163
transform 1 0 9108 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_91
timestamp 1667941163
transform 1 0 9476 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_98
timestamp 1667941163
transform 1 0 10120 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_106
timestamp 1667941163
transform 1 0 10856 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_122
timestamp 1667941163
transform 1 0 12328 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_135
timestamp 1667941163
transform 1 0 13524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_141
timestamp 1667941163
transform 1 0 14076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_151
timestamp 1667941163
transform 1 0 14996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1667941163
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1667941163
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_180
timestamp 1667941163
transform 1 0 17664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_187
timestamp 1667941163
transform 1 0 18308 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_9
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_16
timestamp 1667941163
transform 1 0 2576 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1667941163
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_73
timestamp 1667941163
transform 1 0 7820 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_110
timestamp 1667941163
transform 1 0 11224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_124
timestamp 1667941163
transform 1 0 12512 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1667941163
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_147
timestamp 1667941163
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_151
timestamp 1667941163
transform 1 0 14996 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1667941163
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_181
timestamp 1667941163
transform 1 0 17756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1667941163
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_384
timestamp 1667941163
transform 1 0 36432 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_12
timestamp 1667941163
transform 1 0 2208 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_19
timestamp 1667941163
transform 1 0 2852 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_31
timestamp 1667941163
transform 1 0 3956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_43
timestamp 1667941163
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_82
timestamp 1667941163
transform 1 0 8648 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_94
timestamp 1667941163
transform 1 0 9752 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 1667941163
transform 1 0 10304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_103
timestamp 1667941163
transform 1 0 10580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1667941163
transform 1 0 12512 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_143
timestamp 1667941163
transform 1 0 14260 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1667941163
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_174
timestamp 1667941163
transform 1 0 17112 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_180
timestamp 1667941163
transform 1 0 17664 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_192
timestamp 1667941163
transform 1 0 18768 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_204
timestamp 1667941163
transform 1 0 19872 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1667941163
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_16
timestamp 1667941163
transform 1 0 2576 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_107
timestamp 1667941163
transform 1 0 10948 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_118
timestamp 1667941163
transform 1 0 11960 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_126
timestamp 1667941163
transform 1 0 12696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_145
timestamp 1667941163
transform 1 0 14444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_151
timestamp 1667941163
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_158
timestamp 1667941163
transform 1 0 15640 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_164
timestamp 1667941163
transform 1 0 16192 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_176
timestamp 1667941163
transform 1 0 17296 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1667941163
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_385
timestamp 1667941163
transform 1 0 36524 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_11
timestamp 1667941163
transform 1 0 2116 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_23
timestamp 1667941163
transform 1 0 3220 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_35
timestamp 1667941163
transform 1 0 4324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1667941163
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_119
timestamp 1667941163
transform 1 0 12052 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_131
timestamp 1667941163
transform 1 0 13156 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_143
timestamp 1667941163
transform 1 0 14260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1667941163
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_155
timestamp 1667941163
transform 1 0 15364 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_376
timestamp 1667941163
transform 1 0 35696 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_384
timestamp 1667941163
transform 1 0 36432 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_148
timestamp 1667941163
transform 1 0 14720 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_154
timestamp 1667941163
transform 1 0 15272 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_166
timestamp 1667941163
transform 1 0 16376 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_178
timestamp 1667941163
transform 1 0 17480 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp 1667941163
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_385
timestamp 1667941163
transform 1 0 36524 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_14
timestamp 1667941163
transform 1 0 2392 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_26
timestamp 1667941163
transform 1 0 3496 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_38
timestamp 1667941163
transform 1 0 4600 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 1667941163
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_155
timestamp 1667941163
transform 1 0 15364 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_159
timestamp 1667941163
transform 1 0 15732 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1667941163
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_126
timestamp 1667941163
transform 1 0 12696 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1667941163
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_230
timestamp 1667941163
transform 1 0 22264 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_236
timestamp 1667941163
transform 1 0 22816 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1667941163
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_373
timestamp 1667941163
transform 1 0 35420 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_376
timestamp 1667941163
transform 1 0 35696 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_384
timestamp 1667941163
transform 1 0 36432 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1667941163
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_124
timestamp 1667941163
transform 1 0 12512 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_130
timestamp 1667941163
transform 1 0 13064 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_134
timestamp 1667941163
transform 1 0 13432 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_140
timestamp 1667941163
transform 1 0 13984 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_152
timestamp 1667941163
transform 1 0 15088 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1667941163
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_231
timestamp 1667941163
transform 1 0 22356 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_235
timestamp 1667941163
transform 1 0 22724 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_247
timestamp 1667941163
transform 1 0 23828 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_259
timestamp 1667941163
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1667941163
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_217
timestamp 1667941163
transform 1 0 21068 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_222
timestamp 1667941163
transform 1 0 21528 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_234
timestamp 1667941163
transform 1 0 22632 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1667941163
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_385
timestamp 1667941163
transform 1 0 36524 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_102
timestamp 1667941163
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1667941163
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_7
timestamp 1667941163
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1667941163
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_93
timestamp 1667941163
transform 1 0 9660 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_99
timestamp 1667941163
transform 1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_106
timestamp 1667941163
transform 1 0 10856 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_118
timestamp 1667941163
transform 1 0 11960 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_130
timestamp 1667941163
transform 1 0 13064 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_384
timestamp 1667941163
transform 1 0 36432 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1667941163
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_201
timestamp 1667941163
transform 1 0 19596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_213
timestamp 1667941163
transform 1 0 20700 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_225
timestamp 1667941163
transform 1 0 21804 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_237
timestamp 1667941163
transform 1 0 22908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1667941163
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_258
timestamp 1667941163
transform 1 0 24840 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_264
timestamp 1667941163
transform 1 0 25392 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_276
timestamp 1667941163
transform 1 0 26496 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_288
timestamp 1667941163
transform 1 0 27600 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_300
timestamp 1667941163
transform 1 0 28704 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_373
timestamp 1667941163
transform 1 0 35420 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_376
timestamp 1667941163
transform 1 0 35696 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_384
timestamp 1667941163
transform 1 0 36432 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_385
timestamp 1667941163
transform 1 0 36524 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_381
timestamp 1667941163
transform 1 0 36156 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_384
timestamp 1667941163
transform 1 0 36432 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_7
timestamp 1667941163
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1667941163
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_373
timestamp 1667941163
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_384
timestamp 1667941163
transform 1 0 36432 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_14
timestamp 1667941163
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_273
timestamp 1667941163
transform 1 0 26220 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_279
timestamp 1667941163
transform 1 0 26772 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_285
timestamp 1667941163
transform 1 0 27324 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_297
timestamp 1667941163
transform 1 0 28428 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1667941163
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_373
timestamp 1667941163
transform 1 0 35420 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_376
timestamp 1667941163
transform 1 0 35696 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_384
timestamp 1667941163
transform 1 0 36432 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_21
timestamp 1667941163
transform 1 0 3036 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_24
timestamp 1667941163
transform 1 0 3312 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_36
timestamp 1667941163
transform 1 0 4416 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_48
timestamp 1667941163
transform 1 0 5520 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_118
timestamp 1667941163
transform 1 0 11960 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_130
timestamp 1667941163
transform 1 0 13064 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_140
timestamp 1667941163
transform 1 0 13984 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_152
timestamp 1667941163
transform 1 0 15088 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1667941163
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_292
timestamp 1667941163
transform 1 0 27968 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_298
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_306
timestamp 1667941163
transform 1 0 29256 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_318
timestamp 1667941163
transform 1 0 30360 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_365
timestamp 1667941163
transform 1 0 34684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_368
timestamp 1667941163
transform 1 0 34960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_376
timestamp 1667941163
transform 1 0 35696 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_384
timestamp 1667941163
transform 1 0 36432 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_14
timestamp 1667941163
transform 1 0 2392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_22
timestamp 1667941163
transform 1 0 3128 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_43
timestamp 1667941163
transform 1 0 5060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_48
timestamp 1667941163
transform 1 0 5520 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_70
timestamp 1667941163
transform 1 0 7544 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_91
timestamp 1667941163
transform 1 0 9476 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_99
timestamp 1667941163
transform 1 0 10212 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1667941163
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_119
timestamp 1667941163
transform 1 0 12052 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_131
timestamp 1667941163
transform 1 0 13156 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_146
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1667941163
transform 1 0 26036 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_275
timestamp 1667941163
transform 1 0 26404 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_323
timestamp 1667941163
transform 1 0 30820 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_329
timestamp 1667941163
transform 1 0 31372 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1667941163
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_358
timestamp 1667941163
transform 1 0 34040 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_384
timestamp 1667941163
transform 1 0 36432 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 36892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 36892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 36892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 36892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 36892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 36892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 36892 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 36892 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 36892 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 36892 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 36892 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 36892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 36892 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 36892 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 36892 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 36892 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 36892 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 36892 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 36892 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 36892 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 36892 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 36892 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 36892 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 36892 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 36892 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _236_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 6992 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _237_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 11960 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform -1 0 11224 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 10580 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform -1 0 9476 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform -1 0 6808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform -1 0 10488 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform -1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform -1 0 10580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform -1 0 11040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform -1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform -1 0 10212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _248_
timestamp 1667941163
transform 1 0 9200 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform 1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform -1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform 1 0 10120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 4784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform -1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform -1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform -1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform -1 0 19872 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform -1 0 22632 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform 1 0 14168 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform 1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1667941163
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform -1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform 1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform 1 0 20976 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform 1 0 20056 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform -1 0 23460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform -1 0 17388 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform -1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform -1 0 12144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform 1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1667941163
transform -1 0 13800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform -1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform -1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform 1 0 14720 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform 1 0 9568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform -1 0 15364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform -1 0 16192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 13156 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform -1 0 18308 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform -1 0 18308 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform 1 0 9384 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform -1 0 17112 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform 1 0 18400 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 16836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform 1 0 2760 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform 1 0 9844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform 1 0 12420 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform 1 0 14352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform -1 0 2576 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1667941163
transform 1 0 9200 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1667941163
transform -1 0 8740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1667941163
transform -1 0 3588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1667941163
transform 1 0 2668 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1667941163
transform -1 0 7176 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1667941163
transform 1 0 11040 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1667941163
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1667941163
transform 1 0 10488 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1667941163
transform -1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1667941163
transform -1 0 13800 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1667941163
transform 1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1667941163
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1667941163
transform 1 0 15732 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1667941163
transform 1 0 15088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1667941163
transform -1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1667941163
transform 1 0 10672 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1667941163
transform -1 0 15088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1667941163
transform 1 0 13248 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1667941163
transform -1 0 18676 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1667941163
transform -1 0 16376 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1667941163
transform -1 0 16744 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1667941163
transform 1 0 12604 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1667941163
transform 1 0 11776 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1667941163
transform 1 0 17940 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1667941163
transform 1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1667941163
transform -1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1667941163
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1667941163
transform 1 0 12420 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1667941163
transform 1 0 7360 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1667941163
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1667941163
transform -1 0 21068 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1667941163
transform -1 0 22540 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1667941163
transform 1 0 5152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1667941163
transform 1 0 8004 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1667941163
transform -1 0 17480 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1667941163
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1667941163
transform 1 0 6532 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1667941163
transform -1 0 15640 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1667941163
transform -1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1667941163
transform -1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1667941163
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1667941163
transform -1 0 18032 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1667941163
transform -1 0 16376 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1667941163
transform 1 0 10948 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1667941163
transform -1 0 2392 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1667941163
transform -1 0 14536 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1667941163
transform -1 0 14444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1667941163
transform 1 0 11408 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1667941163
transform -1 0 2300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1667941163
transform 1 0 18216 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1667941163
transform 1 0 15456 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1667941163
transform 1 0 6900 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1667941163
transform -1 0 14628 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1667941163
transform 1 0 16928 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1667941163
transform 1 0 12052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1667941163
transform 1 0 6992 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1667941163
transform 1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1667941163
transform 1 0 19044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1667941163
transform -1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1667941163
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1667941163
transform -1 0 14996 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1667941163
transform 1 0 19872 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1667941163
transform 1 0 8648 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1667941163
transform 1 0 12052 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1667941163
transform 1 0 13524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1667941163
transform 1 0 13340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1667941163
transform -1 0 11224 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1667941163
transform 1 0 11592 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1667941163
transform -1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1667941163
transform 1 0 8372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1667941163
transform 1 0 11684 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1667941163
transform 1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1667941163
transform 1 0 16652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1667941163
transform 1 0 12328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1667941163
transform -1 0 12788 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1667941163
transform 1 0 10488 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1667941163
transform -1 0 15732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1667941163
transform -1 0 15272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1667941163
transform 1 0 11500 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1667941163
transform 1 0 12144 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1667941163
transform -1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp 1667941163
transform 1 0 14444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1667941163
transform 1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1667941163
transform -1 0 15640 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1667941163
transform 1 0 11960 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1667941163
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1667941163
transform 1 0 11316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1667941163
transform -1 0 13800 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1667941163
transform 1 0 16008 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1667941163
transform 1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1667941163
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1667941163
transform -1 0 19320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1667941163
transform 1 0 12144 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1667941163
transform -1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1667941163
transform 1 0 2668 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1667941163
transform 1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1667941163
transform 1 0 3404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1667941163
transform 1 0 28612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1667941163
transform -1 0 26496 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1667941163
transform -1 0 12512 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1667941163
transform -1 0 11960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1667941163
transform -1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1667941163
transform -1 0 20976 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1667941163
transform 1 0 3956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1667941163
transform -1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1667941163
transform -1 0 17112 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1667941163
transform -1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1667941163
transform 1 0 10672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1667941163
transform -1 0 18492 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1667941163
transform -1 0 10856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1667941163
transform -1 0 15916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1667941163
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1667941163
transform -1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1667941163
transform -1 0 2208 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _428_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1667941163
transform -1 0 18308 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform -1 0 26404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1667941163
transform -1 0 22264 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform -1 0 17112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform -1 0 22264 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform 1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform 1 0 4784 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1667941163
transform 1 0 13248 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1667941163
transform -1 0 16468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1667941163
transform -1 0 19688 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1667941163
transform -1 0 16376 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1667941163
transform -1 0 13064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1667941163
transform -1 0 10488 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1667941163
transform 1 0 2760 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1667941163
transform 1 0 19320 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1667941163
transform 1 0 21804 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1667941163
transform -1 0 15732 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _447_
timestamp 1667941163
transform -1 0 22724 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform -1 0 25024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform 1 0 22356 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform -1 0 5060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform 1 0 9936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform 1 0 21252 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1667941163
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform -1 0 7360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _455_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _456_
timestamp 1667941163
transform 1 0 9384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1667941163
transform -1 0 8648 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1667941163
transform -1 0 8648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1667941163
transform -1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1667941163
transform 1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1667941163
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1667941163
transform -1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 1667941163
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp 1667941163
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1667941163
transform -1 0 9476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _467_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1667941163
transform -1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1667941163
transform 1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1667941163
transform -1 0 10120 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 1667941163
transform -1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1667941163
transform -1 0 10672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _473_
timestamp 1667941163
transform -1 0 9384 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1667941163
transform -1 0 10304 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1667941163
transform -1 0 10304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1667941163
transform -1 0 10580 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _477_
timestamp 1667941163
transform -1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _478_
timestamp 1667941163
transform -1 0 11224 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _479_
timestamp 1667941163
transform -1 0 9568 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1667941163
transform -1 0 10948 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _481_
timestamp 1667941163
transform -1 0 10028 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _482_
timestamp 1667941163
transform -1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _483_
timestamp 1667941163
transform -1 0 10304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _484_
timestamp 1667941163
transform -1 0 10488 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _485_
timestamp 1667941163
transform -1 0 10028 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1667941163
transform -1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _487_
timestamp 1667941163
transform -1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 1667941163
transform -1 0 10028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _489_
timestamp 1667941163
transform 1 0 10212 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _490_
timestamp 1667941163
transform -1 0 9660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _491_
timestamp 1667941163
transform -1 0 10396 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1667941163
transform -1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _493_
timestamp 1667941163
transform -1 0 6072 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _494_
timestamp 1667941163
transform -1 0 8648 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _495_
timestamp 1667941163
transform -1 0 10304 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _496_
timestamp 1667941163
transform -1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _497_
timestamp 1667941163
transform -1 0 4784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _498_
timestamp 1667941163
transform -1 0 7268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _499_
timestamp 1667941163
transform 1 0 9292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _500_
timestamp 1667941163
transform -1 0 10488 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _501_
timestamp 1667941163
transform -1 0 6072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 1667941163
transform -1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _503_
timestamp 1667941163
transform -1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _504_
timestamp 1667941163
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 1667941163
transform -1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 1667941163
transform -1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 1667941163
transform -1 0 10120 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _508_
timestamp 1667941163
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _509_
timestamp 1667941163
transform -1 0 8004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _510_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _511_
timestamp 1667941163
transform 1 0 1564 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1667941163
transform -1 0 3496 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _513_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 8648 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _514_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _515_
timestamp 1667941163
transform 1 0 7268 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp 1667941163
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _517_
timestamp 1667941163
transform 1 0 6532 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 1667941163
transform -1 0 6072 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _519_
timestamp 1667941163
transform 1 0 7360 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _520_
timestamp 1667941163
transform 1 0 4416 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _521_
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _522_
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _523_
timestamp 1667941163
transform -1 0 3404 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1667941163
transform -1 0 7452 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _525_
timestamp 1667941163
transform 1 0 6716 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _526_
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _527_
timestamp 1667941163
transform -1 0 3680 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 1667941163
transform 1 0 4232 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _529_
timestamp 1667941163
transform -1 0 3772 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _530_
timestamp 1667941163
transform -1 0 8648 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _531_
timestamp 1667941163
transform 1 0 7268 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _532_
timestamp 1667941163
transform 1 0 7636 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _533_
timestamp 1667941163
transform 1 0 6716 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _534_
timestamp 1667941163
transform -1 0 5980 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _535_
timestamp 1667941163
transform 1 0 4232 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _536_
timestamp 1667941163
transform -1 0 3404 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _537_
timestamp 1667941163
transform 1 0 7268 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _538_
timestamp 1667941163
transform -1 0 8648 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _539_
timestamp 1667941163
transform 1 0 7176 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _540_
timestamp 1667941163
transform 1 0 3956 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _541_
timestamp 1667941163
transform 1 0 2208 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _542_
timestamp 1667941163
transform 1 0 6256 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _543_
timestamp 1667941163
transform -1 0 4968 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _544_
timestamp 1667941163
transform 1 0 6532 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _545_
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _546_
timestamp 1667941163
transform 1 0 1656 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _547_
timestamp 1667941163
transform -1 0 3404 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _548_
timestamp 1667941163
transform -1 0 6072 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _549_
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _550_
timestamp 1667941163
transform 1 0 4692 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _551_
timestamp 1667941163
transform 1 0 4048 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _552_
timestamp 1667941163
transform 1 0 1656 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _553_
timestamp 1667941163
transform -1 0 3496 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _554_
timestamp 1667941163
transform 1 0 4232 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _555_
timestamp 1667941163
transform 1 0 1564 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _556_
timestamp 1667941163
transform -1 0 8648 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _557_
timestamp 1667941163
transform 1 0 6532 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _558_
timestamp 1667941163
transform 1 0 1656 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _559_
timestamp 1667941163
transform 1 0 1656 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _560_
timestamp 1667941163
transform -1 0 3496 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _561_
timestamp 1667941163
transform 1 0 7268 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _562_
timestamp 1667941163
transform -1 0 6072 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _563_
timestamp 1667941163
transform 1 0 3036 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _564_
timestamp 1667941163
transform 1 0 1656 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _565_
timestamp 1667941163
transform 1 0 1564 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _566_
timestamp 1667941163
transform -1 0 3404 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _567_
timestamp 1667941163
transform 1 0 7084 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _568_
timestamp 1667941163
transform 1 0 4232 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _569_
timestamp 1667941163
transform 1 0 3312 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _570_
timestamp 1667941163
transform -1 0 3496 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _571_
timestamp 1667941163
transform 1 0 1656 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _572_
timestamp 1667941163
transform -1 0 5612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _573_
timestamp 1667941163
transform 1 0 7544 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _574_
timestamp 1667941163
transform -1 0 8648 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _575_
timestamp 1667941163
transform 1 0 7268 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _576_
timestamp 1667941163
transform 1 0 5704 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _577_
timestamp 1667941163
transform 1 0 4232 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _578_
timestamp 1667941163
transform -1 0 6072 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _579_
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _580_
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _581_
timestamp 1667941163
transform -1 0 3680 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _594_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 36156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _595_
timestamp 1667941163
transform -1 0 36064 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _596_
timestamp 1667941163
transform -1 0 14720 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _597_
timestamp 1667941163
transform -1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _598_
timestamp 1667941163
transform 1 0 2576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _599_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19228 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _600_
timestamp 1667941163
transform -1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _601_
timestamp 1667941163
transform -1 0 27876 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _602_
timestamp 1667941163
transform -1 0 20240 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _603_
timestamp 1667941163
transform -1 0 36156 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _604_
timestamp 1667941163
transform 1 0 16008 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _605_
timestamp 1667941163
transform 1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _606_
timestamp 1667941163
transform -1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _607_
timestamp 1667941163
transform -1 0 26772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _608_
timestamp 1667941163
transform -1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _609_
timestamp 1667941163
transform 1 0 15824 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _610_
timestamp 1667941163
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _611_
timestamp 1667941163
transform -1 0 20424 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _612_
timestamp 1667941163
transform 1 0 15088 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _613_
timestamp 1667941163
transform 1 0 2300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _614_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _615_
timestamp 1667941163
transform 1 0 10028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _616_
timestamp 1667941163
transform -1 0 18952 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _617_
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _618_
timestamp 1667941163
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _619_
timestamp 1667941163
transform 1 0 4784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _620_
timestamp 1667941163
transform -1 0 19136 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _621_
timestamp 1667941163
transform 1 0 12236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _622_
timestamp 1667941163
transform -1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _623_
timestamp 1667941163
transform 1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _624_
timestamp 1667941163
transform 1 0 14628 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _625_
timestamp 1667941163
transform -1 0 26128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _626_
timestamp 1667941163
transform -1 0 31372 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _627_
timestamp 1667941163
transform -1 0 17204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _628_
timestamp 1667941163
transform -1 0 27416 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _629_
timestamp 1667941163
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _630_
timestamp 1667941163
transform 1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _631_
timestamp 1667941163
transform 1 0 13156 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _632_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 15640 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _633_
timestamp 1667941163
transform 1 0 12328 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _634_
timestamp 1667941163
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _635_
timestamp 1667941163
transform 1 0 12880 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _636_
timestamp 1667941163
transform -1 0 18952 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _636__92 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18768 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _637_
timestamp 1667941163
transform -1 0 20792 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _638_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _639_
timestamp 1667941163
transform 1 0 14260 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _640_
timestamp 1667941163
transform 1 0 12972 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _641_
timestamp 1667941163
transform -1 0 17572 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _642_
timestamp 1667941163
transform 1 0 12788 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _643_
timestamp 1667941163
transform 1 0 13524 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _644_
timestamp 1667941163
transform -1 0 16284 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _645_
timestamp 1667941163
transform 1 0 16744 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _646_
timestamp 1667941163
transform 1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _647_
timestamp 1667941163
transform -1 0 14720 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _648__93
timestamp 1667941163
transform -1 0 17204 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _648_
timestamp 1667941163
transform 1 0 17572 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _649_
timestamp 1667941163
transform 1 0 12972 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _650_
timestamp 1667941163
transform 1 0 11316 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _651_
timestamp 1667941163
transform 1 0 10580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _652_
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _653_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _654_
timestamp 1667941163
transform -1 0 15640 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _655_
timestamp 1667941163
transform -1 0 12604 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _656_
timestamp 1667941163
transform 1 0 13432 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _657_
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _658_
timestamp 1667941163
transform 1 0 5612 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _659__94
timestamp 1667941163
transform 1 0 11684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _659_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _660_
timestamp 1667941163
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _661_
timestamp 1667941163
transform -1 0 15088 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _662_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _663_
timestamp 1667941163
transform -1 0 13800 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _664_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _665_
timestamp 1667941163
transform -1 0 11224 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _666_
timestamp 1667941163
transform 1 0 11684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _667_
timestamp 1667941163
transform 1 0 12052 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _668_
timestamp 1667941163
transform 1 0 16560 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _669_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _670_
timestamp 1667941163
transform 1 0 13984 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _671__95
timestamp 1667941163
transform -1 0 18676 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _671_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _672_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _673_
timestamp 1667941163
transform -1 0 20516 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _674_
timestamp 1667941163
transform 1 0 12420 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _675_
timestamp 1667941163
transform -1 0 17664 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _676_
timestamp 1667941163
transform 1 0 14628 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _677_
timestamp 1667941163
transform 1 0 17572 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _678_
timestamp 1667941163
transform 1 0 14168 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _679_
timestamp 1667941163
transform -1 0 13984 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _680_
timestamp 1667941163
transform -1 0 4140 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _681_
timestamp 1667941163
transform -1 0 2392 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _682_
timestamp 1667941163
transform 1 0 12052 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _683_
timestamp 1667941163
transform 1 0 12604 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _683__96
timestamp 1667941163
transform -1 0 12236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _684_
timestamp 1667941163
transform -1 0 15824 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _685_
timestamp 1667941163
transform -1 0 19964 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _686_
timestamp 1667941163
transform -1 0 11500 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _687_
timestamp 1667941163
transform -1 0 16376 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _688_
timestamp 1667941163
transform -1 0 2668 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _689_
timestamp 1667941163
transform 1 0 14168 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _690_
timestamp 1667941163
transform -1 0 18768 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _691_
timestamp 1667941163
transform -1 0 16192 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _692_
timestamp 1667941163
transform -1 0 13708 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _693_
timestamp 1667941163
transform 1 0 9384 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _694_
timestamp 1667941163
transform -1 0 21252 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _695_
timestamp 1667941163
transform -1 0 16376 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _695__97
timestamp 1667941163
transform -1 0 16008 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _696_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _697_
timestamp 1667941163
transform 1 0 19780 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _698_
timestamp 1667941163
transform -1 0 21344 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _699_
timestamp 1667941163
transform -1 0 21068 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _700_
timestamp 1667941163
transform -1 0 13524 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _701_
timestamp 1667941163
transform 1 0 8740 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _702_
timestamp 1667941163
transform -1 0 15180 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _703_
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _704_
timestamp 1667941163
transform 1 0 16652 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _705_
timestamp 1667941163
transform 1 0 17204 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _706_
timestamp 1667941163
transform -1 0 20700 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _707__98
timestamp 1667941163
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _707_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _708_
timestamp 1667941163
transform 1 0 13064 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _709_
timestamp 1667941163
transform -1 0 16376 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _710_
timestamp 1667941163
transform 1 0 15548 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _711_
timestamp 1667941163
transform 1 0 15272 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _712_
timestamp 1667941163
transform 1 0 17848 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _713_
timestamp 1667941163
transform 1 0 12696 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _714_
timestamp 1667941163
transform -1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _715_
timestamp 1667941163
transform -1 0 18952 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _716_
timestamp 1667941163
transform -1 0 12236 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _717_
timestamp 1667941163
transform -1 0 13248 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _718_
timestamp 1667941163
transform -1 0 16100 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _719_
timestamp 1667941163
transform 1 0 15180 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _719__99
timestamp 1667941163
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _720_
timestamp 1667941163
transform -1 0 13708 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _721_
timestamp 1667941163
transform 1 0 11316 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _722_
timestamp 1667941163
transform -1 0 11224 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _723_
timestamp 1667941163
transform -1 0 13616 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _724_
timestamp 1667941163
transform -1 0 11224 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _725_
timestamp 1667941163
transform -1 0 16284 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _726_
timestamp 1667941163
transform -1 0 15732 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _727_
timestamp 1667941163
transform -1 0 12972 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _728_
timestamp 1667941163
transform 1 0 5244 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _729_
timestamp 1667941163
transform 1 0 5060 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _730_
timestamp 1667941163
transform -1 0 2392 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _731_
timestamp 1667941163
transform 1 0 7820 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _731__100
timestamp 1667941163
transform 1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _732_
timestamp 1667941163
transform 1 0 11868 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _733_
timestamp 1667941163
transform -1 0 13340 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _734_
timestamp 1667941163
transform -1 0 15088 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _735_
timestamp 1667941163
transform -1 0 13800 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _736_
timestamp 1667941163
transform -1 0 8372 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _737_
timestamp 1667941163
transform -1 0 10028 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _738_
timestamp 1667941163
transform 1 0 6808 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _739_
timestamp 1667941163
transform -1 0 10764 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _740_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _741_
timestamp 1667941163
transform 1 0 14996 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _742_
timestamp 1667941163
transform 1 0 14076 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _743_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _743__101
timestamp 1667941163
transform -1 0 16468 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _744_
timestamp 1667941163
transform 1 0 18032 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _745_
timestamp 1667941163
transform -1 0 20240 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _746_
timestamp 1667941163
transform 1 0 11776 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _747_
timestamp 1667941163
transform 1 0 12972 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _748_
timestamp 1667941163
transform 1 0 14352 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _749_
timestamp 1667941163
transform 1 0 17848 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _750_
timestamp 1667941163
transform 1 0 15088 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _751_
timestamp 1667941163
transform -1 0 15088 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _752_
timestamp 1667941163
transform -1 0 12512 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _753_
timestamp 1667941163
transform -1 0 10672 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _754_
timestamp 1667941163
transform -1 0 12236 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _755_
timestamp 1667941163
transform -1 0 13432 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _755__102
timestamp 1667941163
transform -1 0 13064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _756_
timestamp 1667941163
transform 1 0 15364 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _757_
timestamp 1667941163
transform 1 0 19872 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _758_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _759_
timestamp 1667941163
transform -1 0 17388 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _760_
timestamp 1667941163
transform -1 0 11960 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _761_
timestamp 1667941163
transform -1 0 13432 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _762_
timestamp 1667941163
transform -1 0 21988 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _763_
timestamp 1667941163
transform -1 0 16836 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _764_
timestamp 1667941163
transform -1 0 14996 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _765_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _766_
timestamp 1667941163
transform -1 0 21896 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _767__103
timestamp 1667941163
transform 1 0 20700 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _767_
timestamp 1667941163
transform -1 0 20332 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _768_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _769_
timestamp 1667941163
transform 1 0 19872 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _770_
timestamp 1667941163
transform -1 0 20608 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _771_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _772_
timestamp 1667941163
transform -1 0 15088 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _773_
timestamp 1667941163
transform 1 0 11408 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _774_
timestamp 1667941163
transform 1 0 22264 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _775_
timestamp 1667941163
transform -1 0 19688 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4232 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1667941163
transform 1 0 2576 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1667941163
transform 1 0 2576 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1667941163
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1667941163
transform 1 0 4324 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1667941163
transform -1 0 10948 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1667941163
transform -1 0 3496 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1667941163
transform -1 0 6164 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1667941163
transform 1 0 4232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1667941163
transform -1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1667941163
transform -1 0 33304 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform -1 0 36432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1667941163
transform -1 0 36432 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1667941163
transform -1 0 36432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform -1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform -1 0 1840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform -1 0 1840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform -1 0 15272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1667941163
transform -1 0 36432 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1667941163
transform -1 0 36432 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform -1 0 36432 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform -1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform -1 0 35236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1667941163
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform -1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform -1 0 36432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 5244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 36156 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform -1 0 36432 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform -1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform -1 0 36432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1667941163
transform -1 0 36432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform -1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform -1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform -1 0 36432 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform 1 0 36064 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform 1 0 36064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform 1 0 36064 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 3128 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform -1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 36064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform 1 0 36064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform 1 0 23276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform 1 0 35512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform -1 0 13800 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform 1 0 36064 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform -1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform -1 0 1932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 36064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform -1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform -1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform -1 0 10764 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform -1 0 3404 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform -1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 36064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 35328 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 36064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform -1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 2668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 36064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform -1 0 2392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform -1 0 9476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform -1 0 4324 0 1 9792
box -38 -48 406 592
<< labels >>
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
port 0 nsew signal tristate
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
port 1 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
port 2 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
port 3 nsew signal tristate
flabel metal3 s 37200 688 37800 808 0 FreeSans 480 0 0 0 ccff_head
port 4 nsew signal input
flabel metal3 s 37200 14288 37800 14408 0 FreeSans 480 0 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 37200 21088 37800 21208 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 37200 32648 37800 32768 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 37200 27888 37800 28008 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 16 nsew signal input
flabel metal3 s 200 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 17 nsew signal input
flabel metal3 s 37200 34688 37800 34808 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 18 nsew signal input
flabel metal3 s 37200 8848 37800 8968 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 19 nsew signal input
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 20 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 21 nsew signal input
flabel metal3 s 37200 29248 37800 29368 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 22 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 23 nsew signal input
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_left_in[9]
port 24 nsew signal input
flabel metal3 s 37200 5448 37800 5568 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 25 nsew signal tristate
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 26 nsew signal tristate
flabel metal3 s 37200 31288 37800 31408 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 27 nsew signal tristate
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 28 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 29 nsew signal tristate
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 30 nsew signal tristate
flabel metal2 s 7746 200 7802 800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 31 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 32 nsew signal tristate
flabel metal3 s 37200 25848 37800 25968 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 33 nsew signal tristate
flabel metal3 s 37200 10888 37800 11008 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 34 nsew signal tristate
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal3 s 37200 36048 37800 36168 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal3 s 37200 17688 37800 17808 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 44 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 45 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chanx_right_in[11]
port 46 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 47 nsew signal input
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_right_in[13]
port 48 nsew signal input
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chanx_right_in[14]
port 49 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chanx_right_in[15]
port 50 nsew signal input
flabel metal2 s 10966 200 11022 800 0 FreeSans 224 90 0 0 chanx_right_in[16]
port 51 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_right_in[17]
port 52 nsew signal input
flabel metal3 s 37200 15648 37800 15768 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 53 nsew signal input
flabel metal3 s 37200 7488 37800 7608 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 54 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 55 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 56 nsew signal input
flabel metal3 s 37200 2048 37800 2168 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 57 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 58 nsew signal input
flabel metal3 s 37200 12248 37800 12368 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 59 nsew signal input
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 60 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 61 nsew signal input
flabel metal3 s 37200 24488 37800 24608 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 62 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 63 nsew signal tristate
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 chanx_right_out[10]
port 64 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 65 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chanx_right_out[12]
port 66 nsew signal tristate
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 67 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 68 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 69 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 70 nsew signal tristate
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 71 nsew signal tristate
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 72 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal3 s 37200 38088 37800 38208 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal3 s 37200 4088 37800 4208 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 pReset
port 82 nsew signal input
flabel metal3 s 200 14968 800 15088 0 FreeSans 480 0 0 0 prog_clk
port 83 nsew signal input
flabel metal3 s 37200 22448 37800 22568 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
port 84 nsew signal tristate
flabel metal2 s 20626 200 20682 800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_
port 85 nsew signal tristate
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_
port 86 nsew signal tristate
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_
port 87 nsew signal tristate
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_
port 88 nsew signal tristate
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_
port 89 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_
port 90 nsew signal tristate
flabel metal3 s 200 11568 800 11688 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_
port 91 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 vccd1
port 92 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 92 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 92 nsew signal bidirectional
flabel metal3 s 37200 19048 37800 19168 0 FreeSans 480 0 0 0 vssd1
port 93 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 93 nsew signal bidirectional
rlabel metal1 18998 37536 18998 37536 0 vccd1
rlabel metal1 18998 36992 18998 36992 0 vssd1
rlabel metal1 6992 7718 6992 7718 0 _000_
rlabel metal2 8510 9554 8510 9554 0 _001_
rlabel metal1 7774 8534 7774 8534 0 _002_
rlabel metal2 6946 10914 6946 10914 0 _003_
rlabel metal1 10580 12954 10580 12954 0 _004_
rlabel metal2 2898 12988 2898 12988 0 _005_
rlabel metal2 2990 5746 2990 5746 0 _006_
rlabel metal1 5152 5066 5152 5066 0 _007_
rlabel metal1 4462 6426 4462 6426 0 _008_
rlabel metal1 9115 16150 9115 16150 0 _009_
rlabel metal1 6716 17306 6716 17306 0 _010_
rlabel metal1 7176 11866 7176 11866 0 _011_
rlabel metal1 2990 15511 2990 15511 0 _012_
rlabel metal1 2698 18666 2698 18666 0 _013_
rlabel metal1 6916 23018 6916 23018 0 _014_
rlabel metal1 8747 19754 8747 19754 0 _015_
rlabel metal2 9614 22593 9614 22593 0 _016_
rlabel metal2 7498 12019 7498 12019 0 _017_
rlabel metal1 10051 22406 10051 22406 0 _018_
rlabel metal1 3687 18326 3687 18326 0 _019_
rlabel metal2 8004 23324 8004 23324 0 _020_
rlabel metal2 10810 19176 10810 19176 0 _021_
rlabel metal1 9529 22678 9529 22678 0 _022_
rlabel metal1 8977 17578 8977 17578 0 _023_
rlabel metal1 6263 18326 6263 18326 0 _024_
rlabel metal2 9522 20519 9522 20519 0 _025_
rlabel via1 2530 9641 2530 9641 0 _026_
rlabel metal2 9246 15368 9246 15368 0 _027_
rlabel metal2 7866 13367 7866 13367 0 _028_
rlabel metal1 9844 13974 9844 13974 0 _029_
rlabel metal1 8372 18938 8372 18938 0 _030_
rlabel metal1 8234 18054 8234 18054 0 _031_
rlabel metal1 8832 17782 8832 17782 0 _032_
rlabel metal1 4745 16150 4745 16150 0 _033_
rlabel metal1 8372 16558 8372 16558 0 _034_
rlabel metal1 8970 17714 8970 17714 0 _035_
rlabel metal2 2070 8738 2070 8738 0 _036_
rlabel metal2 2622 7038 2622 7038 0 _037_
rlabel metal2 7038 11220 7038 11220 0 _038_
rlabel metal1 9660 9622 9660 9622 0 _039_
rlabel metal1 5842 16082 5842 16082 0 _040_
rlabel metal1 6348 18394 6348 18394 0 _041_
rlabel metal1 6302 9146 6302 9146 0 _042_
rlabel metal1 2744 13226 2744 13226 0 _043_
rlabel metal1 6401 13974 6401 13974 0 _044_
rlabel metal2 9982 13056 9982 13056 0 _045_
rlabel metal1 8057 15402 8057 15402 0 _046_
rlabel metal3 6900 13124 6900 13124 0 _047_
rlabel metal1 4239 14314 4239 14314 0 _048_
rlabel metal1 4055 13974 4055 13974 0 _049_
rlabel via2 2714 19771 2714 19771 0 _050_
rlabel metal2 10442 21080 10442 21080 0 _051_
rlabel metal2 5290 18904 5290 18904 0 _052_
rlabel metal1 5244 15062 5244 15062 0 _053_
rlabel metal1 10304 17306 10304 17306 0 _054_
rlabel metal1 4009 16490 4009 16490 0 _055_
rlabel metal2 8142 13209 8142 13209 0 _056_
rlabel metal1 9161 13974 9161 13974 0 _057_
rlabel metal1 5941 15402 5941 15402 0 _058_
rlabel metal1 8740 21658 8740 21658 0 _059_
rlabel metal2 2070 5542 2070 5542 0 _060_
rlabel metal2 3082 6596 3082 6596 0 _061_
rlabel metal2 5290 7140 5290 7140 0 _062_
rlabel metal2 8510 10472 8510 10472 0 _063_
rlabel metal2 9338 10336 9338 10336 0 _064_
rlabel metal1 10948 15130 10948 15130 0 _065_
rlabel metal1 5980 6358 5980 6358 0 _066_
rlabel metal2 5934 8228 5934 8228 0 _067_
rlabel metal2 5014 7548 5014 7548 0 _068_
rlabel metal1 5796 8602 5796 8602 0 _069_
rlabel metal1 1748 5882 1748 5882 0 _070_
rlabel metal2 2898 12653 2898 12653 0 _071_
rlabel metal1 1794 5712 1794 5712 0 _072_
rlabel metal1 10028 12750 10028 12750 0 _073_
rlabel metal1 6578 17170 6578 17170 0 _074_
rlabel metal1 10212 20910 10212 20910 0 _075_
rlabel metal2 21666 17510 21666 17510 0 _076_
rlabel metal1 10028 12818 10028 12818 0 _077_
rlabel metal1 10488 13294 10488 13294 0 _078_
rlabel metal2 1978 4352 1978 4352 0 _079_
rlabel metal1 15732 16218 15732 16218 0 _080_
rlabel metal2 12282 21896 12282 21896 0 _081_
rlabel metal1 18124 12886 18124 12886 0 _082_
rlabel metal2 12006 17646 12006 17646 0 _083_
rlabel metal2 18722 17170 18722 17170 0 _084_
rlabel metal1 17802 17850 17802 17850 0 _085_
rlabel metal1 12006 16626 12006 16626 0 _086_
rlabel metal2 14398 15096 14398 15096 0 _087_
rlabel metal1 13202 24072 13202 24072 0 _088_
rlabel metal1 17342 13192 17342 13192 0 _089_
rlabel metal1 13386 22406 13386 22406 0 _090_
rlabel metal2 13754 17272 13754 17272 0 _091_
rlabel metal2 14674 10268 14674 10268 0 _092_
rlabel metal2 16974 16354 16974 16354 0 _093_
rlabel metal2 11914 20264 11914 20264 0 _094_
rlabel metal2 15134 20264 15134 20264 0 _095_
rlabel metal1 14950 13430 14950 13430 0 _096_
rlabel metal1 12972 11866 12972 11866 0 _097_
rlabel metal1 11408 22202 11408 22202 0 _098_
rlabel metal1 10718 22066 10718 22066 0 _099_
rlabel metal1 12650 12954 12650 12954 0 _100_
rlabel metal1 17802 10710 17802 10710 0 _101_
rlabel metal2 15410 18904 15410 18904 0 _102_
rlabel metal2 12650 22848 12650 22848 0 _103_
rlabel metal2 13570 24616 13570 24616 0 _104_
rlabel metal1 13110 27064 13110 27064 0 _105_
rlabel metal1 6118 24378 6118 24378 0 _106_
rlabel metal1 11822 26554 11822 26554 0 _107_
rlabel metal1 13202 17544 13202 17544 0 _108_
rlabel metal1 13386 19448 13386 19448 0 _109_
rlabel metal1 13984 23630 13984 23630 0 _110_
rlabel metal1 13616 22066 13616 22066 0 _111_
rlabel metal2 14490 24378 14490 24378 0 _112_
rlabel metal2 10994 26520 10994 26520 0 _113_
rlabel metal1 11868 15130 11868 15130 0 _114_
rlabel metal1 12236 25330 12236 25330 0 _115_
rlabel metal2 16974 25177 16974 25177 0 _116_
rlabel metal1 8050 22746 8050 22746 0 _117_
rlabel metal2 15042 14824 15042 14824 0 _118_
rlabel metal2 19642 23256 19642 23256 0 _119_
rlabel metal1 17020 21658 17020 21658 0 _120_
rlabel metal2 20286 23902 20286 23902 0 _121_
rlabel metal2 12650 19822 12650 19822 0 _122_
rlabel metal2 17066 25704 17066 25704 0 _123_
rlabel metal2 14858 24174 14858 24174 0 _124_
rlabel metal2 17802 25432 17802 25432 0 _125_
rlabel metal1 14628 26214 14628 26214 0 _126_
rlabel metal1 14076 20910 14076 20910 0 _127_
rlabel metal2 3910 24174 3910 24174 0 _128_
rlabel metal1 2208 24378 2208 24378 0 _129_
rlabel metal1 12282 13192 12282 13192 0 _130_
rlabel metal1 13570 16490 13570 16490 0 _131_
rlabel metal2 15594 21352 15594 21352 0 _132_
rlabel metal1 19550 16150 19550 16150 0 _133_
rlabel metal2 11270 25432 11270 25432 0 _134_
rlabel metal1 16192 19482 16192 19482 0 _135_
rlabel metal1 2300 23290 2300 23290 0 _136_
rlabel metal2 14398 12648 14398 12648 0 _137_
rlabel metal2 17342 15912 17342 15912 0 _138_
rlabel metal1 17388 23290 17388 23290 0 _139_
rlabel metal1 12926 26214 12926 26214 0 _140_
rlabel metal1 9614 24072 9614 24072 0 _141_
rlabel metal1 20930 16762 20930 16762 0 _142_
rlabel metal2 16146 23902 16146 23902 0 _143_
rlabel metal2 22218 19550 22218 19550 0 _144_
rlabel metal2 21298 18904 21298 18904 0 _145_
rlabel metal2 22402 17918 22402 17918 0 _146_
rlabel metal1 20884 24378 20884 24378 0 _147_
rlabel metal2 13294 25330 13294 25330 0 _148_
rlabel metal2 8970 24174 8970 24174 0 _149_
rlabel metal2 14950 27166 14950 27166 0 _150_
rlabel metal2 19642 20026 19642 20026 0 _151_
rlabel metal2 16882 9962 16882 9962 0 _152_
rlabel via2 12742 11339 12742 11339 0 _153_
rlabel metal1 19320 15130 19320 15130 0 _154_
rlabel metal1 18032 13498 18032 13498 0 _155_
rlabel metal1 12926 16150 12926 16150 0 _156_
rlabel metal1 16422 12886 16422 12886 0 _157_
rlabel metal1 16652 23290 16652 23290 0 _158_
rlabel metal1 15870 13498 15870 13498 0 _159_
rlabel metal2 18078 11288 18078 11288 0 _160_
rlabel metal2 12926 21182 12926 21182 0 _161_
rlabel via1 17805 12138 17805 12138 0 _162_
rlabel metal1 18630 26282 18630 26282 0 _163_
rlabel metal1 11546 14042 11546 14042 0 _164_
rlabel metal2 13018 12410 13018 12410 0 _165_
rlabel metal2 15870 16728 15870 16728 0 _166_
rlabel metal1 15318 13498 15318 13498 0 _167_
rlabel metal1 14214 19482 14214 19482 0 _168_
rlabel metal1 11546 18632 11546 18632 0 _169_
rlabel metal2 10994 22440 10994 22440 0 _170_
rlabel metal2 13662 14824 13662 14824 0 _171_
rlabel metal1 10810 12410 10810 12410 0 _172_
rlabel metal2 15870 10472 15870 10472 0 _173_
rlabel metal1 15226 11866 15226 11866 0 _174_
rlabel metal1 13294 23834 13294 23834 0 _175_
rlabel metal1 4462 23766 4462 23766 0 _176_
rlabel metal2 5290 26180 5290 26180 0 _177_
rlabel metal2 2254 24344 2254 24344 0 _178_
rlabel metal2 8602 26520 8602 26520 0 _179_
rlabel metal2 12098 18734 12098 18734 0 _180_
rlabel metal2 13110 19176 13110 19176 0 _181_
rlabel metal1 14674 22678 14674 22678 0 _182_
rlabel metal1 13064 22202 13064 22202 0 _183_
rlabel metal1 7498 23766 7498 23766 0 _184_
rlabel metal1 9568 26010 9568 26010 0 _185_
rlabel metal2 7038 24786 7038 24786 0 _186_
rlabel metal2 10534 25262 10534 25262 0 _187_
rlabel metal1 14950 22712 14950 22712 0 _188_
rlabel metal1 15226 22984 15226 22984 0 _189_
rlabel metal1 13984 13498 13984 13498 0 _190_
rlabel metal1 17618 19414 17618 19414 0 _191_
rlabel metal1 17618 21114 17618 21114 0 _192_
rlabel metal1 18952 19482 18952 19482 0 _193_
rlabel metal2 13018 14960 13018 14960 0 _194_
rlabel metal1 15686 14586 15686 14586 0 _195_
rlabel metal1 10442 21046 10442 21046 0 _196_
rlabel metal1 18124 22746 18124 22746 0 _197_
rlabel metal1 16146 18326 16146 18326 0 _198_
rlabel metal2 15226 21250 15226 21250 0 _199_
rlabel metal1 11776 8602 11776 8602 0 _200_
rlabel metal1 9430 7514 9430 7514 0 _201_
rlabel metal2 12006 10200 12006 10200 0 _202_
rlabel metal2 13202 8024 13202 8024 0 _203_
rlabel metal1 15594 15368 15594 15368 0 _204_
rlabel metal1 19734 15062 19734 15062 0 _205_
rlabel metal1 11960 21658 11960 21658 0 _206_
rlabel metal1 17342 20026 17342 20026 0 _207_
rlabel metal1 10948 8058 10948 8058 0 _208_
rlabel metal2 13202 10200 13202 10200 0 _209_
rlabel metal1 21758 18632 21758 18632 0 _210_
rlabel metal1 16928 23154 16928 23154 0 _211_
rlabel metal1 13708 9010 13708 9010 0 _212_
rlabel metal2 14490 11288 14490 11288 0 _213_
rlabel metal1 21758 13498 21758 13498 0 _214_
rlabel metal1 20148 12614 20148 12614 0 _215_
rlabel metal1 22770 13974 22770 13974 0 _216_
rlabel metal1 20148 13498 20148 13498 0 _217_
rlabel metal2 22494 13668 22494 13668 0 _218_
rlabel metal1 17802 13974 17802 13974 0 _219_
rlabel metal1 14076 9146 14076 9146 0 _220_
rlabel metal1 11362 17306 11362 17306 0 _221_
rlabel metal2 22494 14178 22494 14178 0 _222_
rlabel metal1 19596 11866 19596 11866 0 _223_
rlabel metal1 11776 37094 11776 37094 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
rlabel metal1 24656 37094 24656 37094 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
rlabel metal2 4554 1520 4554 1520 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
rlabel metal3 1188 4828 1188 4828 0 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
rlabel metal2 36386 1853 36386 1853 0 ccff_head
rlabel metal2 36294 14297 36294 14297 0 ccff_tail
rlabel metal1 32706 37434 32706 37434 0 chanx_left_in[0]
rlabel metal2 36294 21335 36294 21335 0 chanx_left_in[10]
rlabel metal2 36294 32759 36294 32759 0 chanx_left_in[11]
rlabel via2 1610 32011 1610 32011 0 chanx_left_in[12]
rlabel metal1 14260 2414 14260 2414 0 chanx_left_in[13]
rlabel metal1 18216 37230 18216 37230 0 chanx_left_in[14]
rlabel metal2 36294 27999 36294 27999 0 chanx_left_in[15]
rlabel metal2 36754 1928 36754 1928 0 chanx_left_in[16]
rlabel metal2 1610 28883 1610 28883 0 chanx_left_in[17]
rlabel metal1 1150 36142 1150 36142 0 chanx_left_in[18]
rlabel metal1 14674 37434 14674 37434 0 chanx_left_in[1]
rlabel metal2 4002 5984 4002 5984 0 chanx_left_in[2]
rlabel via2 36386 34731 36386 34731 0 chanx_left_in[3]
rlabel via2 36294 8891 36294 8891 0 chanx_left_in[4]
rlabel metal1 26496 37434 26496 37434 0 chanx_left_in[5]
rlabel metal1 9798 2346 9798 2346 0 chanx_left_in[6]
rlabel metal2 36294 29427 36294 29427 0 chanx_left_in[7]
rlabel metal1 30544 2414 30544 2414 0 chanx_left_in[8]
rlabel metal1 34224 37434 34224 37434 0 chanx_left_in[9]
rlabel via2 36294 5525 36294 5525 0 chanx_left_out[0]
rlabel metal1 21758 37094 21758 37094 0 chanx_left_out[10]
rlabel metal2 35834 31637 35834 31637 0 chanx_left_out[11]
rlabel metal2 2898 37961 2898 37961 0 chanx_left_out[12]
rlabel metal3 1188 1428 1188 1428 0 chanx_left_out[13]
rlabel metal2 1702 17867 1702 17867 0 chanx_left_out[14]
rlabel metal2 7774 1520 7774 1520 0 chanx_left_out[15]
rlabel metal1 16928 37094 16928 37094 0 chanx_left_out[16]
rlabel metal3 36532 25908 36532 25908 0 chanx_left_out[17]
rlabel metal2 36294 11101 36294 11101 0 chanx_left_out[18]
rlabel metal1 23368 37094 23368 37094 0 chanx_left_out[1]
rlabel metal3 1188 3468 1188 3468 0 chanx_left_out[2]
rlabel metal2 35466 1520 35466 1520 0 chanx_left_out[3]
rlabel metal2 13570 38158 13570 38158 0 chanx_left_out[4]
rlabel metal2 36294 36057 36294 36057 0 chanx_left_out[5]
rlabel metal2 23874 1520 23874 1520 0 chanx_left_out[6]
rlabel metal3 1188 20468 1188 20468 0 chanx_left_out[7]
rlabel metal3 1188 27268 1188 27268 0 chanx_left_out[8]
rlabel metal2 36294 17901 36294 17901 0 chanx_left_out[9]
rlabel metal2 1702 37145 1702 37145 0 chanx_right_in[0]
rlabel metal1 32384 2346 32384 2346 0 chanx_right_in[10]
rlabel metal2 16146 1554 16146 1554 0 chanx_right_in[11]
rlabel metal1 27232 2346 27232 2346 0 chanx_right_in[12]
rlabel metal1 36846 36822 36846 36822 0 chanx_right_in[13]
rlabel metal1 5336 37230 5336 37230 0 chanx_right_in[14]
rlabel metal1 3312 2278 3312 2278 0 chanx_right_in[15]
rlabel metal2 11086 2125 11086 2125 0 chanx_right_in[16]
rlabel metal1 33626 2346 33626 2346 0 chanx_right_in[17]
rlabel metal2 36386 15895 36386 15895 0 chanx_right_in[18]
rlabel metal2 36294 7667 36294 7667 0 chanx_right_in[1]
rlabel metal2 2806 5491 2806 5491 0 chanx_right_in[2]
rlabel metal2 1610 35343 1610 35343 0 chanx_right_in[3]
rlabel metal2 35834 2805 35834 2805 0 chanx_right_in[4]
rlabel metal2 7130 38260 7130 38260 0 chanx_right_in[5]
rlabel metal2 35834 12563 35834 12563 0 chanx_right_in[6]
rlabel metal2 1610 23953 1610 23953 0 chanx_right_in[7]
rlabel metal1 29072 2278 29072 2278 0 chanx_right_in[8]
rlabel metal2 36386 24463 36386 24463 0 chanx_right_in[9]
rlabel metal3 1188 30668 1188 30668 0 chanx_right_out[0]
rlabel metal1 4002 37094 4002 37094 0 chanx_right_out[10]
rlabel metal2 19366 1520 19366 1520 0 chanx_right_out[11]
rlabel metal2 46 1656 46 1656 0 chanx_right_out[12]
rlabel metal2 22586 1520 22586 1520 0 chanx_right_out[13]
rlabel metal1 10442 37094 10442 37094 0 chanx_right_out[14]
rlabel metal1 20148 37094 20148 37094 0 chanx_right_out[15]
rlabel metal2 2806 14807 2806 14807 0 chanx_right_out[16]
rlabel metal2 3174 25177 3174 25177 0 chanx_right_out[17]
rlabel metal3 1188 21828 1188 21828 0 chanx_right_out[18]
rlabel metal2 1334 1520 1334 1520 0 chanx_right_out[1]
rlabel metal1 36202 37094 36202 37094 0 chanx_right_out[2]
rlabel metal1 28198 37094 28198 37094 0 chanx_right_out[3]
rlabel metal2 17434 1520 17434 1520 0 chanx_right_out[4]
rlabel metal2 35558 37519 35558 37519 0 chanx_right_out[5]
rlabel metal2 36294 4301 36294 4301 0 chanx_right_out[6]
rlabel metal1 4416 10234 4416 10234 0 chanx_right_out[7]
rlabel metal3 1556 17068 1556 17068 0 chanx_right_out[8]
rlabel metal2 6486 1520 6486 1520 0 chanx_right_out[9]
rlabel metal1 2668 8534 2668 8534 0 clknet_0_prog_clk
rlabel metal2 1702 10268 1702 10268 0 clknet_3_0__leaf_prog_clk
rlabel metal1 1656 11118 1656 11118 0 clknet_3_1__leaf_prog_clk
rlabel metal1 5014 11186 5014 11186 0 clknet_3_2__leaf_prog_clk
rlabel metal1 5658 13396 5658 13396 0 clknet_3_3__leaf_prog_clk
rlabel metal2 1610 16932 1610 16932 0 clknet_3_4__leaf_prog_clk
rlabel metal1 2254 22644 2254 22644 0 clknet_3_5__leaf_prog_clk
rlabel metal1 7406 15980 7406 15980 0 clknet_3_6__leaf_prog_clk
rlabel metal2 5934 19312 5934 19312 0 clknet_3_7__leaf_prog_clk
rlabel metal2 13754 22542 13754 22542 0 mem_bottom_ipin_0.DFFR_0_.Q
rlabel metal1 15318 17748 15318 17748 0 mem_bottom_ipin_0.DFFR_1_.Q
rlabel metal2 6578 11713 6578 11713 0 mem_bottom_ipin_0.DFFR_2_.Q
rlabel metal1 2116 12410 2116 12410 0 mem_bottom_ipin_0.DFFR_3_.Q
rlabel metal1 4508 12886 4508 12886 0 mem_bottom_ipin_0.DFFR_4_.Q
rlabel metal1 9568 16694 9568 16694 0 mem_bottom_ipin_0.DFFR_5_.Q
rlabel metal2 12558 20944 12558 20944 0 mem_bottom_ipin_1.DFFR_0_.Q
rlabel metal1 6946 17510 6946 17510 0 mem_bottom_ipin_1.DFFR_1_.Q
rlabel metal2 12466 9010 12466 9010 0 mem_bottom_ipin_1.DFFR_2_.Q
rlabel metal1 10902 12886 10902 12886 0 mem_bottom_ipin_1.DFFR_3_.Q
rlabel metal1 8326 9656 8326 9656 0 mem_bottom_ipin_1.DFFR_4_.Q
rlabel metal1 3404 15062 3404 15062 0 mem_bottom_ipin_1.DFFR_5_.Q
rlabel metal1 1610 15096 1610 15096 0 mem_bottom_ipin_2.DFFR_0_.Q
rlabel metal1 13248 23698 13248 23698 0 mem_bottom_ipin_2.DFFR_1_.Q
rlabel metal1 11638 19346 11638 19346 0 mem_bottom_ipin_2.DFFR_2_.Q
rlabel metal2 5980 20978 5980 20978 0 mem_bottom_ipin_2.DFFR_3_.Q
rlabel metal1 1518 18938 1518 18938 0 mem_bottom_ipin_2.DFFR_4_.Q
rlabel metal1 5750 24786 5750 24786 0 mem_bottom_ipin_2.DFFR_5_.Q
rlabel metal2 14444 23188 14444 23188 0 mem_bottom_ipin_3.DFFR_0_.Q
rlabel metal1 13478 21352 13478 21352 0 mem_bottom_ipin_3.DFFR_1_.Q
rlabel via1 8326 18683 8326 18683 0 mem_bottom_ipin_3.DFFR_2_.Q
rlabel metal1 6946 18938 6946 18938 0 mem_bottom_ipin_3.DFFR_3_.Q
rlabel metal1 2254 18394 2254 18394 0 mem_bottom_ipin_3.DFFR_4_.Q
rlabel metal1 6440 20026 6440 20026 0 mem_bottom_ipin_3.DFFR_5_.Q
rlabel metal1 17940 23086 17940 23086 0 mem_bottom_ipin_4.DFFR_0_.Q
rlabel metal1 15870 21998 15870 21998 0 mem_bottom_ipin_4.DFFR_1_.Q
rlabel metal1 19596 17578 19596 17578 0 mem_bottom_ipin_4.DFFR_2_.Q
rlabel metal2 2530 22593 2530 22593 0 mem_bottom_ipin_4.DFFR_3_.Q
rlabel metal1 2254 23732 2254 23732 0 mem_bottom_ipin_4.DFFR_4_.Q
rlabel metal1 1932 19278 1932 19278 0 mem_bottom_ipin_4.DFFR_5_.Q
rlabel metal2 15594 24004 15594 24004 0 mem_bottom_ipin_5.DFFR_0_.Q
rlabel metal2 22494 19873 22494 19873 0 mem_bottom_ipin_5.DFFR_1_.Q
rlabel metal1 21298 24038 21298 24038 0 mem_bottom_ipin_5.DFFR_2_.Q
rlabel metal1 8004 22202 8004 22202 0 mem_bottom_ipin_5.DFFR_3_.Q
rlabel metal1 4508 22746 4508 22746 0 mem_bottom_ipin_5.DFFR_4_.Q
rlabel metal1 5382 21862 5382 21862 0 mem_bottom_ipin_5.DFFR_5_.Q
rlabel metal1 20102 16150 20102 16150 0 mem_bottom_ipin_6.DFFR_0_.Q
rlabel metal1 16054 24242 16054 24242 0 mem_bottom_ipin_6.DFFR_1_.Q
rlabel metal1 16330 13328 16330 13328 0 mem_bottom_ipin_6.DFFR_2_.Q
rlabel metal1 13294 11764 13294 11764 0 mem_bottom_ipin_6.DFFR_3_.Q
rlabel metal1 11914 8908 11914 8908 0 mem_bottom_ipin_6.DFFR_4_.Q
rlabel metal1 12535 11118 12535 11118 0 mem_bottom_ipin_6.DFFR_5_.Q
rlabel metal2 14490 17748 14490 17748 0 mem_bottom_ipin_7.DFFR_0_.Q
rlabel metal1 16238 17136 16238 17136 0 mem_bottom_ipin_7.DFFR_1_.Q
rlabel metal1 13662 14382 13662 14382 0 mem_bottom_ipin_7.DFFR_2_.Q
rlabel metal2 6026 13532 6026 13532 0 mem_bottom_ipin_7.DFFR_3_.Q
rlabel metal1 2070 13498 2070 13498 0 mem_bottom_ipin_7.DFFR_4_.Q
rlabel metal1 5106 12614 5106 12614 0 mem_bottom_ipin_7.DFFR_5_.Q
rlabel metal1 5842 18802 5842 18802 0 mem_top_ipin_0.DFFR_0_.Q
rlabel metal1 13294 19720 13294 19720 0 mem_top_ipin_0.DFFR_1_.Q
rlabel metal1 9200 21454 9200 21454 0 mem_top_ipin_0.DFFR_2_.Q
rlabel metal1 2162 20026 2162 20026 0 mem_top_ipin_0.DFFR_3_.Q
rlabel metal1 2392 23630 2392 23630 0 mem_top_ipin_0.DFFR_4_.Q
rlabel metal2 3634 18020 3634 18020 0 mem_top_ipin_0.DFFR_5_.Q
rlabel metal1 18492 22610 18492 22610 0 mem_top_ipin_1.DFFR_0_.Q
rlabel metal1 13248 14382 13248 14382 0 mem_top_ipin_1.DFFR_1_.Q
rlabel metal1 18354 19822 18354 19822 0 mem_top_ipin_1.DFFR_2_.Q
rlabel metal1 1794 16762 1794 16762 0 mem_top_ipin_1.DFFR_3_.Q
rlabel metal2 3358 18564 3358 18564 0 mem_top_ipin_1.DFFR_4_.Q
rlabel via2 3450 20587 3450 20587 0 mem_top_ipin_1.DFFR_5_.Q
rlabel metal2 17342 23834 17342 23834 0 mem_top_ipin_2.DFFR_0_.Q
rlabel metal1 14766 15538 14766 15538 0 mem_top_ipin_2.DFFR_1_.Q
rlabel metal1 17296 19822 17296 19822 0 mem_top_ipin_2.DFFR_2_.Q
rlabel metal2 3818 7650 3818 7650 0 mem_top_ipin_2.DFFR_3_.Q
rlabel metal2 3450 8160 3450 8160 0 mem_top_ipin_2.DFFR_4_.Q
rlabel metal1 3542 12750 3542 12750 0 mem_top_ipin_2.DFFR_5_.Q
rlabel metal1 1978 12750 1978 12750 0 mem_top_ipin_3.DFFR_0_.Q
rlabel metal2 22218 13906 22218 13906 0 mem_top_ipin_3.DFFR_1_.Q
rlabel metal1 20056 13294 20056 13294 0 mem_top_ipin_3.DFFR_2_.Q
rlabel metal2 12558 8857 12558 8857 0 mem_top_ipin_3.DFFR_3_.Q
rlabel metal1 12489 8942 12489 8942 0 mem_top_ipin_3.DFFR_4_.Q
rlabel metal1 12788 24242 12788 24242 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal2 11086 24004 11086 24004 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal1 15272 13838 15272 13838 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel metal1 17894 12308 17894 12308 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal2 3956 22080 3956 22080 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal1 16606 12750 16606 12750 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal2 3542 25568 3542 25568 0 mux_bottom_ipin_0.INVTX1_6_.out
rlabel metal1 20608 15538 20608 15538 0 mux_bottom_ipin_0.INVTX1_7_.out
rlabel metal1 13110 22474 13110 22474 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14260 16014 14260 16014 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 17388 18870 17388 18870 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 28980 22542 28980 22542 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 10626 24922 10626 24922 0 mux_bottom_ipin_1.INVTX1_2_.out
rlabel metal2 19642 22304 19642 22304 0 mux_bottom_ipin_1.INVTX1_3_.out
rlabel metal1 13570 23154 13570 23154 0 mux_bottom_ipin_1.INVTX1_4_.out
rlabel metal2 11822 20128 11822 20128 0 mux_bottom_ipin_1.INVTX1_5_.out
rlabel metal2 16974 9588 16974 9588 0 mux_bottom_ipin_1.INVTX1_6_.out
rlabel metal1 17618 16626 17618 16626 0 mux_bottom_ipin_1.INVTX1_7_.out
rlabel metal2 12236 20026 12236 20026 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14444 18666 14444 18666 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 18078 15572 18078 15572 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 13662 12648 13662 12648 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 13800 21454 13800 21454 0 mux_bottom_ipin_2.INVTX1_2_.out
rlabel via2 2346 5627 2346 5627 0 mux_bottom_ipin_2.INVTX1_3_.out
rlabel metal2 13110 16490 13110 16490 0 mux_bottom_ipin_2.INVTX1_4_.out
rlabel metal2 15226 19006 15226 19006 0 mux_bottom_ipin_2.INVTX1_5_.out
rlabel metal1 10902 26418 10902 26418 0 mux_bottom_ipin_2.INVTX1_6_.out
rlabel metal1 2484 24718 2484 24718 0 mux_bottom_ipin_2.INVTX1_7_.out
rlabel metal1 14260 24106 14260 24106 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 13340 23154 13340 23154 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 8234 25942 8234 25942 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 24610 32844 24610 32844 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 17526 25024 17526 25024 0 mux_bottom_ipin_3.INVTX1_2_.out
rlabel metal1 16790 26758 16790 26758 0 mux_bottom_ipin_3.INVTX1_3_.out
rlabel metal1 17756 23630 17756 23630 0 mux_bottom_ipin_3.INVTX1_4_.out
rlabel metal1 20838 23630 20838 23630 0 mux_bottom_ipin_3.INVTX1_5_.out
rlabel metal1 17940 25330 17940 25330 0 mux_bottom_ipin_3.INVTX1_6_.out
rlabel metal1 14168 14926 14168 14926 0 mux_bottom_ipin_3.INVTX1_7_.out
rlabel metal2 14766 25092 14766 25092 0 mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 18676 23766 18676 23766 0 mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19826 23188 19826 23188 0 mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 17250 24684 17250 24684 0 mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 19550 19924 19550 19924 0 mux_bottom_ipin_4.INVTX1_2_.out
rlabel metal1 18998 16014 18998 16014 0 mux_bottom_ipin_4.INVTX1_3_.out
rlabel metal1 15548 15538 15548 15538 0 mux_bottom_ipin_4.INVTX1_4_.out
rlabel metal1 20056 14926 20056 14926 0 mux_bottom_ipin_4.INVTX1_5_.out
rlabel via1 13846 11322 13846 11322 0 mux_bottom_ipin_4.INVTX1_6_.out
rlabel metal2 12098 10523 12098 10523 0 mux_bottom_ipin_4.INVTX1_7_.out
rlabel metal1 15502 21590 15502 21590 0 mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15042 20808 15042 20808 0 mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 2392 25806 2392 25806 0 mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 2024 25806 2024 25806 0 mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 21758 25330 21758 25330 0 mux_bottom_ipin_5.INVTX1_2_.out
rlabel metal2 15686 28016 15686 28016 0 mux_bottom_ipin_5.INVTX1_3_.out
rlabel metal2 22126 18564 22126 18564 0 mux_bottom_ipin_5.INVTX1_4_.out
rlabel metal1 19734 18054 19734 18054 0 mux_bottom_ipin_5.INVTX1_5_.out
rlabel metal1 11040 17714 11040 17714 0 mux_bottom_ipin_5.INVTX1_6_.out
rlabel metal1 21436 17102 21436 17102 0 mux_bottom_ipin_5.INVTX1_7_.out
rlabel metal1 20378 25432 20378 25432 0 mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 22402 19244 22402 19244 0 mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 17043 23494 17043 23494 0 mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 12742 25058 12742 25058 0 mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 17894 26282 17894 26282 0 mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15962 12716 15962 12716 0 mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 17250 17578 17250 17578 0 mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 18998 11050 18998 11050 0 mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 11224 14926 11224 14926 0 mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 12144 18666 12144 18666 0 mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 15686 15776 15686 15776 0 mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 11454 14348 11454 14348 0 mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 13202 23018 13202 23018 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 12650 18462 12650 18462 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 2231 24650 2231 24650 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 7866 31790 7866 31790 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 14490 21828 14490 21828 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 17480 22542 17480 22542 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 18262 24276 18262 24276 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 19412 22678 19412 22678 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 16008 24106 16008 24106 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16652 15470 16652 15470 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 12581 10166 12581 10166 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 9614 8398 9614 8398 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 19274 13260 19274 13260 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 23046 14280 23046 14280 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 20332 12070 20332 12070 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 14306 9690 14306 9690 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 36202 4794 36202 4794 0 net1
rlabel metal2 1794 26622 1794 26622 0 net10
rlabel metal2 7958 26656 7958 26656 0 net100
rlabel metal1 16698 18802 16698 18802 0 net101
rlabel metal1 13156 6426 13156 6426 0 net102
rlabel metal1 20470 12138 20470 12138 0 net103
rlabel metal1 2162 36278 2162 36278 0 net11
rlabel metal2 15042 31552 15042 31552 0 net12
rlabel metal1 10442 16150 10442 16150 0 net13
rlabel metal1 22494 29614 22494 29614 0 net14
rlabel metal2 36110 9384 36110 9384 0 net15
rlabel metal2 27462 37026 27462 37026 0 net16
rlabel metal1 25806 4114 25806 4114 0 net17
rlabel metal1 36110 29478 36110 29478 0 net18
rlabel via2 22586 16099 22586 16099 0 net19
rlabel metal1 13662 30226 13662 30226 0 net2
rlabel metal2 24702 23698 24702 23698 0 net20
rlabel via3 1909 36244 1909 36244 0 net21
rlabel metal1 22816 14790 22816 14790 0 net22
rlabel metal1 17710 2550 17710 2550 0 net23
rlabel metal2 14490 25143 14490 25143 0 net24
rlabel metal2 36202 36215 36202 36215 0 net25
rlabel metal1 4140 37162 4140 37162 0 net26
rlabel metal1 5773 2618 5773 2618 0 net27
rlabel metal1 14214 28526 14214 28526 0 net28
rlabel metal1 25254 18258 25254 18258 0 net29
rlabel metal2 36202 21046 36202 21046 0 net3
rlabel metal1 36064 15878 36064 15878 0 net30
rlabel metal1 20010 22610 20010 22610 0 net31
rlabel metal2 2438 4964 2438 4964 0 net32
rlabel metal2 2714 31484 2714 31484 0 net33
rlabel metal2 19734 16830 19734 16830 0 net34
rlabel metal1 26496 36142 26496 36142 0 net35
rlabel metal1 22448 6290 22448 6290 0 net36
rlabel metal1 1748 22746 1748 22746 0 net37
rlabel metal2 29854 10778 29854 10778 0 net38
rlabel metal2 35926 23358 35926 23358 0 net39
rlabel metal1 22586 17612 22586 17612 0 net4
rlabel metal2 13018 4998 13018 4998 0 net40
rlabel metal1 11270 37230 11270 37230 0 net41
rlabel metal1 23000 30906 23000 30906 0 net42
rlabel metal1 7406 2346 7406 2346 0 net43
rlabel metal1 1886 5168 1886 5168 0 net44
rlabel metal1 35995 14382 35995 14382 0 net45
rlabel via3 15341 24956 15341 24956 0 net46
rlabel metal1 20194 21896 20194 21896 0 net47
rlabel metal2 27830 27812 27830 27812 0 net48
rlabel metal1 3174 37230 3174 37230 0 net49
rlabel metal1 2346 32334 2346 32334 0 net5
rlabel metal1 2162 3026 2162 3026 0 net50
rlabel metal1 1702 17170 1702 17170 0 net51
rlabel metal1 7682 2822 7682 2822 0 net52
rlabel metal2 16882 32980 16882 32980 0 net53
rlabel metal1 36064 20570 36064 20570 0 net54
rlabel metal2 36110 12138 36110 12138 0 net55
rlabel metal1 23092 37230 23092 37230 0 net56
rlabel metal2 3910 4250 3910 4250 0 net57
rlabel metal2 16054 25024 16054 25024 0 net58
rlabel metal1 13984 36550 13984 36550 0 net59
rlabel metal1 16560 2618 16560 2618 0 net6
rlabel metal1 35995 36142 35995 36142 0 net60
rlabel metal2 24610 4284 24610 4284 0 net61
rlabel metal1 1794 26486 1794 26486 0 net62
rlabel via2 1886 27421 1886 27421 0 net63
rlabel metal2 36110 18700 36110 18700 0 net64
rlabel metal2 13202 30532 13202 30532 0 net65
rlabel metal2 4278 37060 4278 37060 0 net66
rlabel metal1 19274 10438 19274 10438 0 net67
rlabel metal1 2668 2414 2668 2414 0 net68
rlabel metal1 22678 2448 22678 2448 0 net69
rlabel metal2 18170 36924 18170 36924 0 net7
rlabel metal1 11224 36890 11224 36890 0 net70
rlabel metal1 19504 37230 19504 37230 0 net71
rlabel metal2 2714 13923 2714 13923 0 net72
rlabel metal1 3680 24378 3680 24378 0 net73
rlabel metal1 2116 21998 2116 21998 0 net74
rlabel metal1 1886 2448 1886 2448 0 net75
rlabel metal2 35650 36788 35650 36788 0 net76
rlabel metal1 27922 36890 27922 36890 0 net77
rlabel metal1 17342 4998 17342 4998 0 net78
rlabel metal1 33350 36754 33350 36754 0 net79
rlabel metal1 18538 25874 18538 25874 0 net8
rlabel metal2 36110 4250 36110 4250 0 net80
rlabel metal2 14582 10999 14582 10999 0 net81
rlabel metal1 6210 12682 6210 12682 0 net82
rlabel metal1 20102 2516 20102 2516 0 net83
rlabel metal1 32430 22610 32430 22610 0 net84
rlabel metal1 20148 3366 20148 3366 0 net85
rlabel metal1 27876 32810 27876 32810 0 net86
rlabel metal2 29118 37060 29118 37060 0 net87
rlabel metal2 2346 33762 2346 33762 0 net88
rlabel metal1 9890 31450 9890 31450 0 net89
rlabel metal2 35466 6528 35466 6528 0 net9
rlabel metal1 25300 2414 25300 2414 0 net90
rlabel metal1 4600 10030 4600 10030 0 net91
rlabel metal1 18768 18394 18768 18394 0 net92
rlabel metal1 17434 14314 17434 14314 0 net93
rlabel metal2 11822 27166 11822 27166 0 net94
rlabel metal2 19550 23392 19550 23392 0 net95
rlabel metal1 12581 16490 12581 16490 0 net96
rlabel metal1 16100 22746 16100 22746 0 net97
rlabel metal1 16882 15062 16882 15062 0 net98
rlabel metal2 14490 14654 14490 14654 0 net99
rlabel metal1 13064 2414 13064 2414 0 pReset
rlabel metal1 4186 14994 4186 14994 0 prog_clk
rlabel via2 36294 22491 36294 22491 0 top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 20654 1520 20654 1520 0 top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 31096 37094 31096 37094 0 top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 29808 37094 29808 37094 0 top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 2070 37094 2070 37094 0 top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_
rlabel metal1 8832 37094 8832 37094 0 top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_
rlabel metal2 25806 1520 25806 1520 0 top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_
rlabel metal1 3956 10166 3956 10166 0 top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_
<< properties >>
string FIXED_BBOX 0 0 38000 40000
<< end >>
